module pslhdsa

import encoding.hex

// The test material parly taken from the test vectors
fn test_slhdsa_internal_signature_verify() ! {
	parameterset := 'SLH-DSA-SHAKE-256s'
	// "signatureinterface": "internal",
	// "tcid": 491
	testpassed := true
	// deferred: false
	sk := '971D294199CE58CAD31A929B27E9EB59CFC3651560128AA5ABDDE2C2C4F39FD67B6943136AFA1F8444638D197781976834507E9D5CBF8EED4F7A8107D471E271A93B0F86E74F2C7FE47EA6A8A9319A074B36BED20D3A9A71D7C8EFF333EE7A6C9455B9F5274810025F02BFC48509DA41C84825011259A29E737291710312BCB8'
	pk := 'A93B0F86E74F2C7FE47EA6A8A9319A074B36BED20D3A9A71D7C8EFF333EE7A6C9455B9F5274810025F02BFC48509DA41C84825011259A29E737291710312BCB8'
	additionalrandomness := '127658FE6BBFADD4DC2A7AC86FB57F044F35573BD1C59BDC35AA61A84805E6BF'
	message := 'E2DF680E1AEB52283252452A9C78F31940BCC7B93F36837A8573E9BEE7DF272155164163CEBFC016EF97715540204F1E69498870273BD6244336CDDB0242BFA3A8854BEB975C62C82CEEF5165AC6B1534EEB00A783D0A6A002D8C03087EC05E4ADCC1CF1739D0A6AF00B40CDDCD8FD036755C707266C6FC477BF89A2C752D36CBCD1EE57CA18A816F32713F3951E5F8B7B87835B59C1B59B23E60A1CB3FD9104FED5EC3C64788AEAB021C8DC0893AB81DB3C9F5856D242A80D53CF54035837BB031C87409F3BC81ADFDA2D9B69C2EFF33B0D75EBB9942085168B772D926AC5DEBD329FF887E78E502859ED77585833848062BFC836F4EEA2140E282D8BF073CC5186F49D477055FAD5ACDFA83734943EB9021E06361664B1D0E668DDE263FC070124ABEC97ED879F69F6DF9BA6BF897CEB0A9187F875F1FD738C8BCE0FBEF0B4478667C0B080494B8A167B2814D73E5BB5779CD318438E68E45C6CE13811B5E41EF372E51A3EF487DDAACB86DED559E06DC3E0C5A30FA7B96B82FEA50727F5559D59FD6DB7AC1F953C3FE2C0FDF9EBE30174082D67523E1C6029913AD331C7C06AC880C9B95B5476F14717E22B08E3FCBCD2D6CFE75F1E1D23B7C80C2310DC54220DC9E0F6A7B6D844F08D857062D32936B44AB086E9CD33A97671703399677ECD8844FE3219B106835CB9B593C7949428FCA58A8FAADD660CFBFAA7AE3A34FEA6204D04F6FB25DB3FD95B6350D92FA31E20AA68970D9F1A8D3BFA58F5F0E0DEBF0A8FC26AB2B4D3643D982FC46AA20654EF988F19F40835E3B8B7ABCE8A19D7081FCDF3E08392B7AFC45CA04283D244E7C9E20FC8E9FE8DFD7046FD6A6497C1DEDBB297AF89D037FE6178178206A529B52210664BF7B2BBB67D7CB1BA911828DBDFA6E8AD8766F72F2E067BA4B40A7921008E838C72A084C35F1E1680006505DC1DCC8D80C72A44A59CD9EC7C761AD593FDB22096F546A86C26AFD7CC0C94091A83F2BF8A9E77D4212578D21B0CAB7337EB2215098089CEDD572BF79B4C691E6FF4F828EA52C0B612BCA11FC423FF981D4B24352A04FD13ABDC124B548A90C3453DF61AA4C9BE5C214C19079434ABF0A280812B0FAF5B660F9DF1A9AEE1032BC336546F14A1189F7633E5856A0DB19D85C12C57B553F99AAC0ABCBD68358F06D2841446D130B1CFD8377F09490871CC5B5ADE3EE7D6B0'
	// hashalg := 'none'
	signature := 'E232E876CDD4006E47B0075067332054DF0EE126DDAB993699AAE83DE87CCCF148B15984CF0531B705073A80ADA871816416A7CC8B692382FEBEC982B99C1847C114BDE38D1953624078148473C29C4ADF36634A0F6ED90CCCDFD9F59DF6941BF10B5034DB242109BC5536626525958A59CBE85E940FC43E1DEFA17AAC3701B9A84E38FE196B081D66C592E0990426D6618BCD3F1969D073C9E27991301AA72D9158D27F585296351CC0B5294C53AE2976034D79F725750730A06F51E91A2D93D22AA622E56B3B276BCF40AF97A59BFA5EE20A6AD63DBA724BFDDB5D85F70331AB9752B8880E7194E45792206ACE81F7FBE3E04049906A35E821613CB8E6263DFEF4BF9D9127632C814451381CF0ACF430DC75FEE5DB41C8D51F3F12AF628E804DE43F7BE0F90100412DAED0C3E8DEBBAD4A549FF171338AA908EC0F4BAFCBA500EAB3082B0505FEF9BC01FC23EC695EA9B538118CAB1B2EACB471F2ED3ECD487D495369CF96B8402EF9F3359F6A65BCFB170F05B2A79968DA4BDA7CC0CAE672D8E8C30F4E1403C87164C89F865A58BCD2E930C158AABE7843B16ED10922E9484669AD5A66B6C62B7C7B4E593ED3D735E3508B01FE9B7F75FC9D489DE979766E09E2677A11D632D323547FD397844C0793FC2594C4A2138DA10E50773FE761B992BEF381A71BB6F8F41E22D6A533B546EBC93245AA6C4CBC01CE2AC341B5D74D653DEF4F1052F92996434B0473BC5963DC98756D93E7E0BB0CEB4DC9599554EBE916CCE32464C2E10D9C5187923F9E4A15B1FED3DEBF2E8FE051C64BC2779B83B0D66AEF1962D6872E4DCD7534CBABF4AA6483205F7DC08157010989751410B8B2E8E08CEF3EC3EA1B15A238A5D2B0E336EB329AD99F8E84CEAED2755BD99547FFE5D780A2B21FB45DDB1943B75875E52BD664F1C5A7B64176C59B881034F630D8BE0C1956604F072A9F9F75152C4704E64AC2193510955576C44EEBD5170A6B6302A08A2217D6CA84DCBB90BF2D00F0756A7662E020150CDF58CE440E0886FCA2AE73313BFD735FAC92B5833157CA49C57B761A7A94F73E2DFFE82FEF5F2EF66A0757C3B9BE8CF0B4E7E013106A1C7A43DD090A1B81B983701AEBEF86AAFB96D6BE0ABDB4E238A680642230748CCFEAA7BE6A81816B7FEB94303E418EB1E22C8ED1965D439122BE873A5E9FC339C0EFC3FFDB694AA16285E1FED0B1C23006D90097D95398D4F347F2090558E047841D56B604AA4213E39B2307C3112877548465116A37590C6ADD12DD68287DC3C04A4E19A9BBCD0228330268C8019BB56523019CEA8B99F6809A7DD8B16300481B2C57CFABF9D9629FA9842995423D54A093C1B0C0F872ABA7EB4E69BA522BA8A5E172F23C82ECD597904054E01C55E47540C5485887CE636465A8A0D33A9AEDD439930D9BDBEDE1CB429E4E9B720684E89252A15A4CDAB78E369268D4CCA07EFEC5A5EB00E1F5F3B134F0AE0D10D91EFB92814AD5D9F2541BFD8073DEF4014C3015FFCEB0E6262912D9C5F0D836B0AE2A0C3E52ACAFAF4E243411D1EE5DB68115651C03074CFD97839EE6E77EA2267FDFE881CE19977C3D2ADBB4C37354A7DA8C0D233391E34AC3B275C3901423F809821C6E98BCD6D9A7009F1CDC1AC1E61C0E60D18B126139627FA0312143F5AB8B2D86991BFD7F9ACD9B0A911393D0B488CE560DAA647D254CEC446CD14FA195A5DC21A796D1DAFDA6BA8A726E2C3A17963EAF13DDC86C8F0912878983EA7509FB2B106940BB4612F1E75C78FB3F86BED54C1939F51097069DA236E3D9E054D7394F99D2A54A900DFE2275818860EB09C175D6FA02C5899F141912BF42F0735FE8EBF53C92BD6FB8E2DEF1A6A85E8F004B0DFC187332869EDF4657106B9379C5FF8B81DBC546C40DA7A0FC8AA48832E37D6A40EB96F012F15983D7A00E90571B1AEDAB74F1679A3BBE57CF4F8F6CF17222875B8B375A9B25C490E8F2E2372FFEB932D1C043F8AAEE96347C4B4C5D046876F30C1436D0F9F9858C12B98DD09254010A3A4B3EDDCA59E2811CFDC4B2692898540D124E710B6F5F315836314213CF88A4703A9949663CD4E16A9E924F0A0964E6621A503B7EC4981517F9C9652FC2FF2D35BE0A6F9CE7D6D258603D3E30B94FBC2B3D37FB8206B3DAAB5F04E0503BAE4F400DC3CAA7348CE442A235ED2ED35971F25E19C237C634F2A23BD6DD187B8FDDAD4B094A6340AFD3E25204E03FA85B3A4815F66D0992A162E35AD016191DEC86D9B1DF42217FF115CB00CD5C99C93D41F26720752690EE4E2329170F23F43F8093C235126573705C59D7107042B0BA3C177EBC347059E838B557B46E7B220849A99D606685D9FE812FEA2613FF15D3935D01381B86E9665772460B2458A39186125E4ED21E9D2C57D59369383D6E47AA05775059AF4FA5EBDF152B02995FF0FB3C04583A8253A4636F1AF0FAD240EB7D005308B84CE45447C40B378F4B0800DA53721661FD9802E3F2BBB02C1DDE9ACF77114DE1A728B5C3FB02A9632CE8B3C32CEE5C57FE2950F5A547D282C5A8F45C529CC01329D5CD634A9EFADCEF68AA306B7D0C203F8486F923EDFE24944BFA55C76466944DF36688DA9816DF32BEEC5053E0D7F6070236187616D363EA27FD92F94B73EE8552CBE28F50DF289A43E43D58B3C5FFBA1B986B615BF6865044745C03E243A7869D285CF6397C38D0EC06AC44AE6349AEDDF657244D5D838D67A78192658D89A7C4DB365D518A9537B42D128D165CD5D811246B7C623E2A2260CA08AED7CE32F09408D7C1D5E43D22439921502175BC02559F516E2BE42C8B1A7B20E0D81A61B43C6CAD7B8823344081791F490B0D4E52B405CEB5D4E3AA9BAA275921094F3E53357FE6E7BC0D4AA09820A55FD75BE0235E374EB3CB69101C3F1583DB076FCAC0C9AE7416816F1540CF2252F67D4A33E0B0C4C6F9AB3C27707665EEDB6F8DA87E0A6F7C9A848C7E6CC65CC378A9B580787EDFDD0971BF7F3739A10A2AB91A6132A736ABF2C88578267E061650193EDA6DD1BC2F3FC32F7489BBCAAADFAD14E282A72EF80A7AD03C604D17C270301F39435A8A3918FE8EBA20342C1FFDC19EFCBBF6F83AA180C30273C4B4474AE1128D45F272FDE0D2A04F2EAA6EFE110D583DCD6867A89E1A12101039056C5630CC6A757AACC01829EF0CB2EE9A813D1DD25EE13F32762EE1EBAC7331DB6ECF896C87FA9AF8A5F992B81FE2A045A142F77AC9C276CBDAA5F5279BDAF8972EBD7D39F244C20D82E8B7555DB57F667C75A488D645103777F4267561D7082AB8C758E745F3A641B9DD84DF5C095F24939EEFE29F11BF30554D1BA4C54B5E9B9B6798709C05200E76C6749C843DFEA67D9F0B73717A2A92C1D7920A5FEEAE093347B0CABEC9717E62A0CF19E1A08F8B8CE1BA2D032652757F07A420C399831D9831677810D3004B143B363FA1981FDFC5512A359C507C3D6322D6FD7A079172F37D5F9FB94B78CFBBA6FCCA8C11504209E691E43B3BD4C1ACD188FCE671ED4EC4B1B09722D175E636CA29FFC84383F61418F63E95E333E83052E01E1BFACFBC173F72A155C694E6A45CFACD691791861070AF72A448165ACA754F0515CA0407671D098D7D9DEB7ACB6361A16A52AFD70259949DAE889F1BAE826C0A5ACA9A875DC5A01B62665415687F40A4882D87F1B30D6C8A84E0536DCDA12AD0606FD56D93E164EE3D52229808E85134787D65291F12DCE86E15315CB65C05B489C079C74B9E62AA661A933D8E44C790F0FD61954079579EB3E71EA6DDC183FA3722E8068321001EE42E4F801309CAA6307D90C2C05C2A4F8D11AF5D4CF62E9244B4CC8B66A86E5BB1A5B198036E9F45DB25C9F1B588443D4ECF8624672335F05DA884A5B5577D16A924DE4CCEE993EFB79D18CD4D48EE715AAFE18797EFB555034DF5808FEE0F59C1B1AE52C017CE4C665FB25B58F0181293E349D172458B8172892F796EC5F00C4CA6137146AA8CEE56318DA39B12F7BE73D25789BC55B02C95FB56172931CFB36A4CF82D604E3A66A86C87C1336DE75EE1ADF1EE71C27DAF549FF975F4A3E0673EF4111C1F253A83D86718F979C6AB01F107A48D0AFC32A7A9BEF8C1BAFA9736A9FD9A8E82326469CFC34AFA6921156366826DAB87540FEC0256EA0135E524EEA55E840EF378DA4B75B33571768AF7A34E95051674DDEF08C8F863961D1C4517F10545EA9515A0C2BA9FC5DEEE86D289DC6F44B7EFAEA9F83F8688699D3718A27FB38FF22324CAC491EB866FD92DD55946B3053A096E248EC3C46F604B3B47A9BED36C49951718EB9C4F286E81BAECEF18C19D44DEA90CECDED89F0C220B7F7000BE0CEDD1B1990A693B4E28EF36F1B34A8A0DEB7C8110F9EAE1A183E4397B55328B118852AC3CBFD92AFFFF3D5FD7F09EA348F48432591E0412BF2ED19D91B2D62070C2E9D8FC3CA0FA8DAD3055CB4351153313A6E8BD05CB0830762C6CB6435D84600308AD1387A7C651913903F10B5058033F04138D38CB1F659855EBFFF992157049A5F107F3B48B4CC26959BCE9E2CF595566D8B666AF8CE7298AECB3F1DDDBBE034D6827E05C7FFD46D42AB53C6C56B68F56EE42A208744C0EC314D645EED7238C35EA437804179C434917AE62D532EC833BB2843C8C389697E797BA26A0CE286E2BA34D0E53B914A3B220F5A8B6A7E0FE2189AD726772884762190D321F59701F951754E031154AA512F759C10BBBB046D86BC71448053349D35E1B49906EB7DA52AC9FF66E08A85BABE186864710CF0EF2168814DBAD297521A2EDE408F76D8901F3493C72127544D7AFE03B2C2B51F6DC97D5A8D35A73F8BC6C13B1EAD25BE3C81FEC7CD79D63DD1FD47911A552FADCD865B92DDE878B72767B2FE65F55DE64F393B3FE1DD906553395395773781F3FD9A6F1420A878848FD4105EF69A666BD85E41C858782115CD96E6550FB96FC9ABECF6E94E77A5CCDF8DA0F7FDD25312DFAC157DEC6BFC3717E0774A97AC36573F5868E06766A023B26F3F6D0D5F35B9A659BA1C79987B61F390B1EFCF24DD2FA331AB09BA46EABA008AA254028441964BA0B76F680FB94774D864D08773BE82980A944A944B46F239F3DBB0CD9F1635301C5AA0998C7C66539173810015D8AA65C5B156E6609345846190B42DF5BE8732D2D6268271C35D678BBECFCFF2FDAAAD1941DFF63781114562BB24A3E5E3A399BC5169BE71E4FEBE78132CBA757046CD5A273812FCB4D9554E6495EF12722AC3BE266DF047C58825F883ACCFA4C30283F0A5DC963FAC460678502D2ABC0344D79666F257AA6233E7AC6F067F03B534FDB2991F65D5FC1D5C0F5222778DCAC6B3A607A0531B7962195F25D128B2E93CEA7D6A03FFA8DE3585F6F83EDB6D1BAB7CFE4600FB8A17E9A0F7C9C17F52D2D53C75FD76C431D42749CA23FD52050D2183D5C29C8AC76605C15031A48B606F484443AB017C2C9221BC91691AD4A2993F49DFC2A8CC61001BE5EE4A7E20FCF07806802196EC25A6F8312D5A9795FC59D8BF25B66C022F38616F696924B9B48871A3314CE2947FB2C47702B090A31A4EFD5EBF180FDB8AD809C42A194C2CAEBC03E28BEC4E580A2810500253CF824F8FD19A3430EB8BC04BB42DE1E30F6FB1038C774E618E0967B6CF0EDE098452564D00C535B33898F16C1F490C60A5F997F98E572276DBC1E9F0DB3B87C5A400F7BAB4158CA4203BEF1E3780717C402E9BD08D5FF45D4E4F6D688539F1DFB53084F3A7EBA757025E4FD27EB75922FE88D137CB1CB70FFAFEB3D3F1671B7A01264087A82F1B470A314FC774E180B20F77750CD9A561786D97F5F35B5AC0C749CA023A1C685E8B9022E369FF866732D6CC56B8270C9865EB3D9035BABAEF3190A23157A62332C2AA95A305AEF83949C999A2D24E6AC1AEBA499F9CEF5BCB18BD0FBD9D5EE52B961AD7E9C8E6AE7AFAE78FF5E1EAC093C1A3FB3F346E9D65546DD8D520699336A54EEF1464FD3267C5B328A2D8BDBC567B2517E43CEBE10879D07A8CBAFA12BFA511E794F1F6F6A9690FFA8AA7969BD42C0F81E263C4C8700575AC068329B57E71627837D15E02A57B23CEE4DC62719F134905680339BFC3AC01197A109855A6223EABE6EA471725458B8F43545AA8F66032383E2783E2B822D2B3EBB16B9559840228BDC9D20CBD67965216D224C66F5B35368D6DE0C66405999CE8A0950B37E10634A13CD1EFF846464CC5FDBF4CF11393168F769D6CB9B0593C43C667D91C9029E514814FDACB44C5DFF9C1C9F79F1381851631451337BE4830E07F9A4B81823FB56071AFF57F0EE08C7C6B02DF1EB2910780575F2BDB9040A1BE68F5B6032CF8943FF129FA53FFD94251277A7F2C1857E19E9EF7488D2CFE99EF95C1FC4892AED7FB5555307F94971F268F2A7327D9A53C6AC90678CA000D4339A0097EC688E5865554A5B0825D8C9D1FFD5B9DEE4C4BC06DEAF4F084C83232D623A78AE39E5DBFB6F2AA5B175B55F3E1BBC6DA85E801F2BB88BE8B39EC7AF8CD725035CDE02865FE4DFD82DD0E7F1843D57297A84EFEFFF08654BE8C2B9184775BBE753138F9C95CA5374D533234F75F57F274D29C96B6E0A83F679BD4F472111E3CF4BF42FB5BA41A4D1BDEA700CFEA9091BD7E04648448C6E5D08CBE7BB2A148BA15A23B7511CD8CAFC6FEED56A673F24D78FCEE6868ABADD916B3862C2B58EA1EB8C0D02456B9FF8FF9A050B9E04B186E6B2C8A823368FB6BA6132474DC47C66A542A411FA9667CA790773D9BBE04830C255D33D687403C0483462F2031E80C51B18978A777C6C7324272DD7F1E814304E6F8E58AF3CC8F4B746B56535AA1B5F62A5E28D0778EF5EC756227BA99C5E30BE8742DAE542E7B837B54A38FB50EA2C006275DB2AD855D2DF56A2FD8B92786018571D5A57736E2A298B6A72082821AD5E7380619AD9166264BD24EFFCA7A0B5807A16EB8CF46879412279F8F5F78909E5CF2D46C232C113E1996BA5BA022A95217172B4FE0A53083D901CC8EA351551625C7FB6258DD57C7E14DE269DF3E96D1B1D6A7E5BE2C991653CC736F362A103885CE506326544336B22E77927F5CFB8924DFB174E82C616374252FFA0C01B4CD1CCF3BEB29FC1AA7A8E643D64D70EAFC715BA22692683418C827CE7D5969E19F125D8EF300536BE43094CBF79E8F249C721C2E8A8486AC77319E4E8D2B37453D873865CF5F60C1BB0746EC8DCB6FAAB59BDE79CA3C18C6C73776F2EA37DD3BB0EE750ECFEB5D950DCAF952892F7E0CA786A326E46A424DF501A68F998903476787146983C72D7498BD12ACDC8F28BC79A0281CE4EE5ADA46208B2B9AA85E7F33019F94FA813A7F2DEAC459D58F6CE31F72C852836B7E4769856389C9C465A2FBA6F0DAD76878FA62D556DFAE78C94DB522BF32AF831D536951EBE7BD00347AAA60D76053474FC33170B5E96F5FDB9C782E7779F9323B7D226FB695649D10D1514CD3498940AF3EE891029DCB22F4768E15CDA56376622EA9055E2F885C91EDC7998D99149CD8B4063CF6A772CFD210E746461AC0E133D6C867410A32F9EAD42B7ECFEDB39665EF14FA02798A727822B854C7F4537C9F9F60988806F3C40D04AB53C9FD96F2C4508CBCF95010A69F5B3E82498D38E226B1C1A69B9E936EA733937A70AECA3B3561A06E998D1A13EFB9920F24A390C8643AA7AE3787A19B331AAE212A2246D79EFEDE29825EEF25CC9D2A20AAE1EBB58683876B522E74C79F2EFDDC791AD9DCAE2251B7AD874A5CA2ACAEC13E403ECF0C664A2C78062B798FEF55BB06CF88C412AB3A5C8917E82F1D0FB2BCCF90F6BCCBF89FD42FA0FA1EA64569852F4265BA3B3EB3FFF2B9AF3F694712DD887FFF010888CDCE65B05B4FD98542372B37B428746F53803AB732BF82052FC836D77B60E2C4650F92D30852DCD45E942FFCCAF638BF6B3D06598FD7D66DCE4947BF7A257DF4D98CFA3219E79E1D665E08208F628F3F36BA4DECB40A6BE65AC3B5EB9656F1DF51EDA5AB285DE17AD93B747F7289237358E94712107BE14DC3512967097AD0871361F0FACA888CB9B066341AA9552F0634625BBF1827BD9D0986C6A2DBC6B6DECBCEA729E1B6C3D6710ACAF110E40FD1E096B1E5ED76D99D6952C977B724BEEFDEBB335602AD442BE35D51F5C7E628294937376502287031B51585053169E1DDD6B46077A5283B411566E88F6AE7AF9D7FB43D693AE705CAFB80CFF77DA6806D8E22950A6EEB70295A3516DB6D61A3A7FF87650FB3EBFC23F8B301CD37AD3709B741DE9D90F915C9D78BB1076601A6F7AB584030CB572FC7B9798071DF57D4916595F884714CAF4A1002FBF0DAF27DCB228D0F87CF9924E092072B2B38307AB4D6E3AD17928EEF83CA255F51FF28CA6E4F59462C2D6354B3BEF124555AE15CA25353BDCB56AA111E987603D461653396FC309A24F11EEF8AA8E04E5548C8FF076A0C20EB88D251903D884B503878AEC07F828F4C9FC8C592EC80F2FD50F33AEB98D26589F93220484959798AC6C2036451F720CECA677C74EA478D89E3B0C7FF4728410F6FD9BE02D32719310A73657F5290A5AC8FBB27BCA9EDB961BDAADABA3AEC27FD34B1464906688BA1059C59C6D6D75A5C59A9FACF4FF927C9814D30014024508433F67345D1FABB17CF274A64BADE21359186DCE4C73806763171032BE5A9F94B28FB470EF4BED3F3ACBFE0C0C174831E4A747DC63FAEBDA6CECAB43DEE8DFA1CB145C4D40B64B2AD66967FF84E45DA5EFB46DCA7253FDBB725B735AA5E1931D16D623B615D7BD298E20EC7FB4A45316B65FA6B85AA41CF9B383D234FE13FD6097EB711E42E4D6C56A204345EEBFC894E62716D53E75E81CFAEC0F6CE20B5C1E9AE2702EDAC7E051C88E91604A07B06663C54125ED4117C2B7B8EB13F9344F6DE4F72BF2FC60689A81513B9786D1679F188E9B75DB2F2B7134698AF2859B405FA083CD5B914111FD5C513CD55D40ADDE71E156B30991829B7CDDBEA5135FD565A2576CBA16738B973C76679D5E090CD6F0C2B8BF801CA57ADE57E06FAE27895C4421C282EB22D46DDEDED8EF93E6D07F864139E13A08EE2E43FEF90123CBB46D2B051D9470350BF057C51FFD541A7674706C58A3A9E99CD6F30F0EDAF1E94F9E442E677DAB829D5540B1A1DF49EFEC880D1A4A37E8D550CC10BE32840C112CCF3E2A62C2CCCF79C391EB4DEB61960E44D3F65C09C093E70C403181F2087F826575F0020039FB4736052BEF4B724C702DE9C6627D7AAC11E6BEDF2711488706280B310716098792803BB0BD9AD59DE40BF46A6DACDFB3E02A1890BA60CCE2ECCB444ED05D08FEB7027A6C893285C7DC95F668926D77DFAC47FD38402AA9AD8BBA9E3B6736381FFB71C7143D0962000C36436FE8763B43BD435A6092F9826D0A6B613D3DF483F1403C4D3AB4388DBBE80397A96F9F4D3A9BA0D706223C843FF9D20B22D1AA9CB1DCF86A09DB2BF68E72183F6E5B2394A723A5A6222CE0166B0A995DE1E869DE574FC0F0053F233F9BC74780B829A7D6BF98941AE5D174DDC0501157D0A4F8415C97B17C8695ABF95AF84BA1BEB6E574BB4B9629AF7FCDF00C74D4B01C1283FBDD83C9C1510B1D50425CE2AFDF2A2B2FB2382C23B4777F669F0E859742B3CFAAD067902626ABE716258A9C155CC3F6E936B7B464F4BC048DCB5AE7488C4951EDB4C439F45489E0ABE1AA577034218024E931CA654C710175CA7E84D887BAEF59B6DDAA7396D53C55B9AB470D37C57970D9FFECBE8E76C86DC3ADB5C28825728C11363EBCACBB40B98EA33163A981A54FAD70718792D88562C9F5AA530FD3602C5730D8D66EF80858F8010C0C4F888086F7FB52A54072034199F648B34824A8EA73F84DB0FCE1DFD85178C86AB03EDDAA11971AA3E6313C0C830FF8AB3AE4979BF047544ABE207C4F15CAF5A2F075E9B72BA6F07C56579637055435FDE7B810A6103A52A061DC4EE4105A432F61FBCAC50C8542E53DFF2AE2786F24B042271658FFCE11441CF6D153B04AB9C1B55027376D4ABD527A4FB30FD58A7EC94C32C7BD761EF16A4F05B2FD2FCF9ECA57F93171222627932B9F6EA33905EB39BA79A946768EF79961BEA8C76A8DF987A9AE7823B87DAAA0EBB47C8B8EB1C94F53112A412282E38555E20234C1891C8D3CB0C32B4DAD843A33D0A0E14B9C00EA2045B1F8BB42A9904862327405BB10D01F13877D6C9E51D27EE1595E4BCE9C5823AB1931967AEF9D6A7E412FAC67B6649AF61556E17CBB974AD26A1135569ADBF0DAA02AF59404FF86963B348031D1A56C05C1F22297685263F26DCF19431C2DE03B84E76BDB23B7060AA13CFD601D2D4543A3FFAA6E70E75A7E6E5FCEE082474F638E68F144AAF94386421C0AD600F5735C5E5F7A42431207925E2533F219B3402CE23DA51FF43A7C5FF786EC9678CE82BC0D9FF819A86CD9222BFF3599C52D328F012F9A7A3F2CBC9FA5AFE46B9FD34758C9C27444CCBEF20839A3B42B449E75BF7E3E4B80E8234A3F76B146AA1FA6D3E9FD3A91C9D527A04EDCAA3BD0A289148CDD720A5139A2C2E08FAD784D260608540F4BE946620C5C9365C81DD0F130F82A7944AB1D322C42612DB2F467AB1C11B3ABC028A34B871FBA5CEED656885A124CAEB500A4DED8776ADBDC2C6CDDAE7AE7BF9B447B76A2C454586C11ABC94DBBCF2FE4038F06504D0BF6E9BE83A2B2B47DDBA8789F974AA61B2697069FC23CF05D27ABF6B03ED9B67646A6AABDE3B46E2223FC3EDC548B62EB2F6AF699C4F564162024DEB7EC84A2E4C303B4A5B044F716D7D374E329F2960EE92E503EFEEA550A4C1C80408CC8E477FD6163AFBE7E0633B18B922E47B21F69169F1C5436BB1C0C76A934AB6A146DB0BB2654AA6EC883A7FEAE2C036D9109BC865F49C0DB0C892FC20CA83496C9A0BB7BF5766D0658A0D79E6B14B033C44C104E52FDF9253F9BFB856EB5A7BEC2B3D7BEAB28368AF2C7AC2ECA8DE3EE1EB24C0758D8334399517C6E0AFD8C3113C04BE12191A8F730C36ABCAFF9BD843987563620A8F7120F7B904D81FE5F49B580A9147A3748A8A4D33C1BB43DCF2E021B0D44574D7F48E791633BEEDD44A932C6A25D803BB393FD7EDD59FC4536FA70EE2E23BACC54856086A56C97E037E0E24196AD3868A4DF92DE0BF92C28ED53B8E2187025289D629F273CF8A58BCAF86C278F0D2776912C293B2108FABA0621DDE3606D21EB635B5ACC41D73EF28A9276F431781AFCD2F1574057328FE8CD747B0C1C9ABD1D8D0EA6BD5AFEB837F185ED9434C823D9B8794CB43DBE5EAF937E7D9C173D1D71BAE41810B9D8DF2759286580912DB081C03E800BC1B2DA7AD7B929C61DE5F949AE7743819C6367DF980F9FC7C2B267F6275A892B54935360669B42B74AC623701D2EEE2955F52A1A62A0FA30E73577375C78A12B050AFF692DD95694864606BC81F8ABFF27B5A7C3A79B05D21A67615EA2185B20B3051D5F70DAD3A3934E80576D35797F3C681865BB3A0A4B3269A1CE147DE6AB0513371BC8C327BAB4793F1DC86AFBEA5C1AEDE5B8B5845D9B1C939430AC8D2E0353353B8C384EE825776A4B15D15595738972287E6EC97593F87E6E6D5485A1FC2C364A3ECD95DDC64258B58092AD4900DD2A0A224F0B2E84AD5AF1FAE5E8D577E9214B16E6FD515F885FD08ACE369F63F8F20198C6860A7B9AC476C42D361F18165B8BD2975972A066C350D89E3E60055D525D3501C3B60C367D9BF3125CD653FEE0CB9217652B920FF9044CB46290AD27A451D5717E21B485A0F1632728A0372BFCB9E43F8E9EAACB48A277B054EB54BADE92A7ABEC5D03293C593D87E71FB90571426CFCF29B80135C518FBFB8686E5F596FADB202531EC239F0D58D7FF2DFF6952FDFB6B5D0DFEFF5717F34CE29614B8E8E08877C4BC87279CCC37088B9F871A16C0A22AC156D70FA386A5AEDF88FD743DEC57CD6CF5531D6B1EB4617663C0E9F8EBD93C22AF81D388053F0C58D6CB09672DB1B72147B228227669A65EF369190F7C35FE0C581EA7EAF68104C6CF8EEAA3949A929FBACFE3EC94A051846457A00FDD8D372364F576262E3D983C9ABA61130FFF11D2AAFEB186F67C58BE01E17A56D302E436E030EB4BE406E7714C55DF94899BC34559D6E4B2A1ACECE1CA3DC021A30551F3F852EE048632A5447731383C00CAA6E880CDF0E5F0E5AC1178BEAC0F25A91B54A476BAE61A549CAA6632E14CADCA9037CE0794527DB3D759722FF0D8B67E05A89D4F1B54B74A68E543BF0E15C5BFC5D7648CCBBD33353F7C5F86A7F47BAE737C6F6F34C10885C0532C89FD37C7D027A758C16BB33F683360668F44D8856A3E56BA277BA4E3E2B180D41B3C68BCCE2563F0E99D38074ED36BEF1C570BB47C7DFC735495F7C39DFAC1B11CDADDA8743AF2613EA4F342F5E8850F7F67AF94224F06659035A102094DB0754BCDE609B24F51BFDD4E9BCF23C922A173CC51215820AA19979D13A5353C1726C5FE6A1D0D7D441D825C31723025BD3AEF60C6B216E7919302ED7A306B4521C20705C6B328BF7563D44C1015CFC2255803ED6D52F2C22691D39F84876099CF3C2CBB6E2568C0EE4DD578FD3E0170885EFA0C2876C1CEA9E46085BF7D0D537E6411FF9F69FEA57622AB85C58F0C1DCF6F3525E1CC32F40C2573D762E61AF007BAA81929B2FAD02F5D7F27AAD8ABA47E114B60F3B491B8B78255DC2A6DBB70FA4F395F94C3CCC977C4F9E7B161BC6FC78DFDA303E7DBC8E749346F5439DF5038551565D0437D81C7A2D8C3E38CDC0666206AD972036AC1511AEB47F23000DDB8C6172C0CC64830C672D13F0D6314837EA04508C4F1D895C8B0B30500D72B486042F7BBBDFC9AA7C63338014305DBFD506189047E61969CD8A1742CFECA9D6F0FFDE9E15E0E25B5B51315FB5090A19A885D10B3FFF9A279F613D20CA496D21BF8952109C30AC226628241371F46AA5875D90D300B2A0AF9B78A8958C18AFB0B037A26CA9062C1B669897AD11409C66BA7469C465D19B5B2759420B5C9F590FDDB0CE5B9DC0B4D14F21B6DE1917EED666E30F587DEF77505F0A3ADEABC18A262BA0CB5D2C022A948E019F40FECA645DB983C153DB3791F654ECD032597927B4D7BEB118A53DC7ED2194163878FC793DE1A4E95F2CFE7C816ED17C2A11E01D2D3EB7C1CC7B895875818C823A579747E1BD48DC3BF895FF566FF98A6E483DFDCE08BE815E2DB540176C0632ABBF0F41D75428F64CFB6AB5BF6B27A6FA6987FEC81D0F48CC0A9FF16876808F3E6EC0779E292B48D5A705F8D07869F17098CE0D83C68E7C15514B589A2E8AAF3ABE6DC42724E359611BC5A10316AD999CB9BF4659B8CEDF96D7501B886D4404E9DCA9C94EC27E08066963ACDA541CB45593BC48073452373D4E5D6AA2330B0200D29EDB9060EC38F9B4AD70F3E52D586BD69832D5BAC7B98995506CAB99CF40B0ED083A6A011D0030AB5D0D1705C23257538FB684C020894CF4D6E1F398EB037C543845B7650CF4C9F356FB5E3BBC9B04D150C797D7699D72F95D0F58036CC6FA8D842A1CE83FFED1E65083C34F066FCD15DABE4AD0A07B8D5B7B7C23FA6F2202149B296C18616E5D902EA625B6E9745293A73511E4D0C979A383B0D611C19237BC1307DAC978CC6DDBA36ACE1CA439FDF140D1A21CC32C3C2DE0785E98EBE706759E164D7E73816EAB53567B348D00368DF3499E5C8B803FF1E986EE489B15B64ABAC894245094786D6EDE852A19C58319134E09B34ABE73D128BA90272964BB4FFFB62ED25F3BE25C38A4EB3362D76CD4E667BA00E2969E73BC4F689DF7FA920016A29E2990BB748F76F04CC86B3333ECB1C4F035CA38F0EDBE7C7E03E94C6645569739B5E3ECA40F9D6120ABB6273B7FC1168C48794F3DFC68E9CA30C9EDF5C7C02109A832029F4A67BB8F2AF1C5C168CF2F6CA91895EA634D44E4D53D82B4F3D1FAD403A6C19EC4CCAACED9D1C98063ED64D657E30B0E9A6AA2D3FC4BAAF6FA078FFFDF2258A69B8843F70A5450C9E256C6DEE4153C4FDE809375FFB60AF02FCBFC4F1BE03349D5730B87CEE5EE1023A85C1858BFAC8D3237527676269E11DBF69898A365BE83B07BFDB4A054B0813C2A385BF628332F9221712F1EAE199C46F2F89C5744F53C8D826C61FD132C40651C04F05FE1C3D2F8867C4B60712E65B523F2FC2134268B93759578DA54B9F6E0B9F083F6BDC32C975F6FAA25A5B61E466A2C5996674730D9C4C12CA7FAB836A4E243A813381E68CD1E37929D25C5C010F8A021BDDA9964609171316389FE915D97B93FEA13437A7A52F5CD38AEF0A33B5502B505B780A32BA3C12817679A84C2B37C58421BE89CB8E0E615E74A23F1738A179FD66F1A34C50DE677A20063A4360F67FD6F8C8854F1E64997BB362C5168896B67AFAA7128E3E3B72A77BE560BB20D0BA7B5E25BEB62E7549784B5E1DAE615646AD301C1EB173FD862DBADB1B49BFBDE3CE944A24747B7BD2CA76DE9488BB9115BAA8B58B64C842AD21235A7AD0666C18B64C7EF9B5FCFAE74F7E0D736517E74C6E976E2394B1DB3FB7FDE5B3157DF933BAF51B45D7D9A23EDE70870BF1F74795705AB2FB31F5C4C00ECD3FCD5D7B12119288802FE04C6671795D2BD24D1D90E63E8766850882BBB17CC0F68311C1C840D0590872C26DA7646785AEE7D3B1044B4D18297F79748F72013D66F1422BA9FFA354408E8A76FCC4569149C9B440A3F695654C484292A3F1AD85A4C6249F47CA4FCF59F2B018D5E5B2D65D738779BD80C4EDDE117A1E62A93D531ABE4DADF2A357D8CA04307C8F0D297645809971B355B325AEDB94BDF305C87B3F3CA4225130914187C6FEBD910201DF6B930233384B9AA29CFFF84A3572FC75AD3D3370ECD23E0D9D000C2D055D69ED81ACBDFB4075C14315DB5519B14C594A9BB01E4AFE56C7AB07D0003999E3F85A69F6719BEF81AAE4BDCB48893E8520300EA36ACDAD079C6F4A03089D77BBFF37DB80167FA973139AEB89514F8B1D002305EC32C051390C895233FB186E343446C7B273AEBA6CADA0A88E57C08575E04EC332462D4530410D90F3AF276D99F9DEB94B6EEFD254E46E6C3009E94150C2AA4D61D21223539B985A0CBAE0025B21955317EA0C1DFC14030FA0A6B3E024DC41AD70B9EDC51EA43C673A3379826AFD852E7E019CEE6788959B0806EE698E307791A9714F07499668CCE4DE6A88FCDC87A90CA5933548087BC02EE559CCF7C55BB63F3AA80D54D0733F202610D81DEE75F1DD1D3C3B776B85311944B79CBA04EAB7993DF3664A71F1DEC2A8BA082EBB3FA2FD4B8339107DD9F15359B8040C55040C5387CB553D7AB7FE31D6EACE1B91B3F7A8B603CDE4C167770D0D4F99E1B43409716F3330B65A6009237772FDB8E8A4A5FED824B7DA15BC8032F36CFD0ABB8C4E7B4156946454D145A23ED16480B40641C71DF650D4A75CB791F9A6BB6E86068D95D62F2AA924C112DADDD68DCD964B7F324A649838068EC8F0E0FD93B55DB1564AF8F7EB862C501471CCA1A5A83F3EDDD7D37F4618B4A6E19CB07D078D049BE6B60526E839F80C5690CC608C1C01F2E24C768EE3E20BD956A6830F95AA08065CC6423E31D29203C669C24F3E209AAC03EC4EDF3843806E3C463ABEEAA22EB476DB63F980D1D0BFA43B372DAE9DF572088E45EC2956F10A346EF000AB5A033C273A6F75FADC1DD9FC8B59B8C56BC3421E13D09325240CCD15AA556E36AB5CD04302CD5E66F350DF4043D09EFD4986AA5B552A63C29FEB41282E1F154CA695E3012563063249002CC34B229449E676A9639FA050A9F2CFF96EFEA88BD38369F81D1366C4842E7655788D11A9D252AABA7616270661E593B64A116825FD73EE2B92DFB9A540FC54D7399597FB46875E7D2BCBC5ABB868CE376C98D55F95F4743A91C852ED559357A2872C72DE1AF3CDE2FA7342C9362924A48BC5071E52F6731BBA7C9EA2289401DC9A1AFE207CD9D81B61024E6C828E2ECA6F6FBB13F84A6BA3B2FDF2D2F59A22AF7B3C21DE80A199CF56B108E08568F8F3004AEC06B2F08533190AE5F4D08BF780FFBB4BFE0840D739E0660692AA174BD39D03A4D7F5D3EE891CC47A306CE286409CD562D96573F74D77A1446CA512FB1D36BC8CDB9927E89BE8AEFCF118C7E613B03B189B303C94CC097C54E28B9D9E6BD3A010DE469A35C18EED4CC063FF3104DCDE1A433E38DA20AF048DB76BF2D63D54D96136C0DADBDAA9FA3ED0C9CD619EB5088A3F947DFD536C8268270474481E4FC7A0AF1AA126262F679F14A914A5B69FACFBC30C8A9E2C86EBB6066A1D24A2A703DBE7599B84919DAFF20E60F9D9B0814F519E56D2FE2806CE532DFF095C2CC93FB989AE58F26D72285EA41E0DA1ABF06FC93A5451C0D153BF46F15B1EF205919673BDCBDC650CDD50EAA79116BA2B2C5ABBF4678A2FFB79F739F0FB508545B395A543AF33652A9C6F0189ABC0AFE966B961D934382B285F39A3BC6630AA2FFE0A9EDC5FA3C2AF1706421280A42AFC91224E6D1EBE43105A9D1D5A6BC97CA38FDB91623A2E332C993C3F127D116CF3ECCFD57BBE0EAAC9A4DD724829B0655861B383A43600180696AC4FDD4724CA385526DA90F7D403AC32EBA82482776392DEE835B95D16ABA7286A87817AF8735916A35439DE1C0EEE7C441A3436D9060547EB09BFDF0158BE66147D9F1526808000E1E9D45613A4A6B3026EFE362F2A1923888F722DDB0F67E6233A86BAC669FB6A9C7C851A1732FB36F14689E9160396BAB78E084584A30578963DA8D78D6ADD68690EB29AB1E6E3A558ADC6219C37A055816024A42AD9F6E5BC897B23D196F016B6B75ACEEA25EE02D0BD3DD36A3A36CEABA9CF766B8A48AB4CB18FB8745EB95C686953FBE590D6E2545CCBA069048502C6148A9C17A25420E4677DBCE37D1B1AAE14E14D6997F6599FF17215306A5446CADEC8291FAF6D20CFE8A05C216C3A2E0BB19143B5C70F274B5E5AB1BD544321E6F1F3780EA31857077A83DA5B0E2BF48E44BEAFFE6D17F86182A49A131EF7F1D3BFF2BFCD00DD09CDBF4AF998E3067A9D17E2CA6FFB7F22F5AFA2F8447CEAAEF938829F99A95FBBECBEB9DD4455A648FD28B3249A86B81896FD760A529291CC2CAEF0B5683A4DE65E9C5EA7B4A3BD5087D141F48A9653568A4830C92DE5ABA7DB492A2E951778B67815D7B6222A65FEA234237D092122E078090DB79190878372B4704F397DD872C5CE5740D8EEF552F92A73A59E9C939A2A6C913966C39D8D9650E782697ED4E40D7F12DCAA550CE1FB2279748FE7D265D9CE800DA696670EAF335B508C2DB3D768E04CEE82162482CD6720C53D3BBB8E61B279FFC0F436B23CDD924A745DA55E773EA28686C3A5DE5B03B2D7BEC3D303CA68D243740EAF3290E309C60C950337BFE39A4CA6B479847993D9427FF025C9DAD84DE6064907E0C1F021F39F5F3BB0EB83A0112FB518173DC287D31B9248E487621F9DB17A64B679445A15AB5C92AFCF622AC37E4EB149A6C7374DB9E4D64F2CC19A4623296732DA95070D1FDA7C8B00FACA6DCD575EE90ECBE73919FE66EDE70C0374CF3117ED3022AE6AF4FD122AA891F23BE99F36AE6269DFB4C4BFAF86B04BD24DF39B07B575984536B809F0EA5EBC1FA5DBFB3C66BD468EB189660538F568DCBAFF11C138C3A91072CFE2A183FD4C75DC698BE7AC8CAE2F8EDD6A821145AA2D0613838AD25F273DC31F0E6C8B7AD66EDB76D715A334BC866FEE4481FDF8900DB2CFEEE7C19249AAF9AECCDD1FEFC55C624E5C8FD67611126B9BFDAF0A7FFDDE12510EBA62A885DB5704484C18D2BB903152E399B4CB48E38B32FA1AFE67FF8411AE69926C770D5603F307BD3B65730F30B936CBBE2564FDC4BCA1947E47B09A7D6A9ACA6CFF14697648C3E2A4CEB1CEE9022ABA62A2034D5CA79AED108AB0824A795E80F881928F1EE686B77B3FB8EB870B607606FA11106BB778012A585E1D08065BBE7040876EDC25759D5E095F8015D57414E7E20A901FB2E685FFA76B04D096C52982F1B22EDF28E8AC648F3E699B9ACEB158305BB5A500C37574E6E4BD760DC1D7F94EA3090430E1B44E61B5FC0F66AABAEDA66BBE44EB371730A4820399EDDC285B7512D8498B4F05DE766D33C64E9D412A1EE532D7E0B5686DBAFBE648F8963839C64A6DBFCB53C271AA89C2E88F91A62491EE65A1DAEFA43CD0EBFC26354077DC4AEB5BFE1C3FD7FFEDD4285847F0AC5F836B4BBD2D3FE8C8B8B67F514AEF14953AFF5E9F74D8C67B6A5EFED7D830DA3910ED427DBDAC890CED62BAA1B3D6AA47AFB498F4AEAAA6A5F84F2626C7FB84FAAE6E96531C89D552A0E105F8A731ABA18AA13A49406E144297FAB457CD5971A5A39778D9EB272409937E7E56936806E4D998AA4E21E76E33262FC4A97D7A2474903AB6794C0B94AB9C0DB350C5E1B320E16C597F22021BC1F937A202B0379A6BBAFC554F6FFCA7CAED3A58F4B5EF727083894216EC9B08849B62D9C1544F4CFCFCA2B7EBD9AF09FB8BB91E0C08AA9C5C6474059ADBFD710EE49673853AD8C84DBBE561FDE5D2EA100B37FFA1D708509957DA52814419095169617EB10B0D4677D567F3D76087B89BABB97F31826F91DA07CE4AFDB4058B3112336F63E6993F8D273DA175783CDDEAAE71426AAC94764BD33A2BA5E54C9266A1596ECDB0062F070B4F2135D916DFE127715EF6E8692829548C799DA25A8C3916CE044654B827F3CF499ADDD3E0850227C9882C565FDCD65E7CBE667840DC64724A6F008B025404B04FDCDFFC6112843717096C06A2970F6E0805B4BCB447C4A9A3A776EA00C4727FDC827766DFB6383869F73B9B393626F48E61FC25C98637F1B46D75EBAFB309C823EB844D7C888ED82D7F2DEB73D485E41F3CF173FE6A27BCD03F442047A7A091D88F3DA2C8819359A3B12D0AF4FAD05279C4C595673E04AA2FFC68EDC9A39DCF7ABF3B57B8C0837C723962369227C96D14F31BE628ADB1779C581D0973B7BD27BBED306C2C35C0AA197C7568847666DD76202B13207625CB96DFFADC203F0A947E320E8C93F20BB015B5A4B5CF625A5B723B1DBE48E5DF7A3821C789DA0343869F24CDA75B0585FC4B5AC626BAF5AB813F5E72AFEA8F9B677B3E0B0527E4B30A085F5B380C29466C88F0B54EC03BC652AB9A9194B12ADC639A3BB40B3CAC6BEC76C17A5A84F2DF084C8EB2F471B5CDD20CDB36448DA3F57615EC7A847CB90414B59E90CF78ED2A4AF09AC520340C1B9DD81FE0D1D8F0E0A0B15D9682FC1B2AD74C0EE461304959E23E86126B0C0F6C0A4A80FAE5896530AEE8D2B22735F3B92716DE54FDAF68355247CF09C694945C9BDC584C9601A9F8427180A64B71EB8803BEF1B0C5A1ED6B23EF585DB9D2A7BE765CA1B48B2FF7758426489A3223B74CF71FA6E6C157BA278E13E408DE2919089C0F588A787B8DF37B2537364E08A6F16D87E65D006B2BD2F2E1C6A94B71777B9132AAFC745B9AE5C1EF173403DCFE6ABADFFE2BDDF6242E935E5D1901EA8B66C228CC21A1DB6BDEFDA845FCE1D52E37538869A7F02BFF0CC2A0ABB544CDAE888B4CE0A6F7B38A5F4D9C559862C01F61F30C4B0D52BDDCDE976710D28F9C38D48A617D8A87BE979CE0CF83181E3A0646BE26F4B6E54C3343A97C12B60A6AC6245743CB40DC1664B421C9A79E83A963D25D1D9C2E9EA4A7D440B2C4253142F8C465447020CDFF391E7F6CFCB860EEC0F207C739194BE4F999B3EE08018D303D7570A82DD3FDE98A4D6700CA49E8F507672406BBDDEDFB7325B2B4CDCA5F5BED2166E3A5C2C377AD25540964DA337157E457A94611906917124C40DFC206ED973ADEC2DD837D0029B8F5B023E527873F6E2603D0208BE75BDEFAF8BAC07D15DD434C40D35AF7B0F2DAC261231ECC9046CBD0333AAA90980B75BC3208FCBE546B03B80B9BE4F46EC6CC5DD4ECB30D49BB05ECAD870DF7E4BA6D890D06E377F848B17E5E26FD1DEF93B0880F1941C486612D4708FDD29B39C5D6E6DED0B23790C2AC963A34946B2E34C2E56494C6B85041B3805F58A20042D7F74FA9E6243084382832EB6D9899D259A191337638EC1BA73FF40A01849D6E748E4EC10218EEEE19A0D99E79370235B554171AF632A9F37A8AEEAE6497C14622D7C43AC458E18A418B0FCB509EED230CAEDFD9F8F2295A63C2B1A93D27577EDEC648EC44E774218D48EEA004E0481E09A09B53C4617FF3B295144544E91D97C38C3AAF098A7B30AD8A4FAE0140052A82A4470B9415FDB4A8077202D7E8BC75F081630A560DA2A60F578DF7B2DFC4923F828D2A469D78172C2974793DFAB8F5DCAABA544B6EDA1D93A7A9BBF8A6E3AAA5688C3E51465DB20FFB2FDAC06095A2855F4FE558B85E44F67C01A8CA44EE6CDB7B0275F823FA600B53E10FAA3C9E4303F53024473848F19E25D013AA529B82FBC90DF4ACF0A36B68EB70890797FE7D4626B95E7C1C27B1E4CD94D8614E197123A3944BEE9D7D7CD336AE8CDF54E4C59219F148B41C479492930B9BD30F53056FA6894A75FCD40404D6C3CD9356BBD09845B4640ABEB828F8952B1D9CE7C0FF0C9A56EF417D782FE5A5FA4D807A001092016CCD4C6AF7A07F64EB3F078DA4A87B906EE0BE3A9C53792F7D4A305CF56524E5FFFE86E3A3211818DF04E30CFAD3DF1B0B09DBED50FB7F731D3A31A192E79A490A36A7E7F323BF90A4235FFE24A8A33A1BAAB8E731479D86DF3D0A0217F1863EDEA243BA5137358119628EF5B1C3B988CD132135781D4D3D90DE8A873A6CF68F9621E6532D336A9F71C9630C9FE22509A74993DC3BFBC792E6BF7D1EB3229FC68C548501E9433AABF1AB544F640E95DC25CBA6AF0BDDD02D37746F7BF72B4AD3417DC17F90CDD341CEE0D036A7A49091A4CA0B71D8F3CAE1BB1CF9C2CBA8E3A3005975A8F5A1AE25D34EC926EC850EB8259C685BCA944D5D000905356352FF2A7BFE636E01E6B7E109A8A2024AD99777015117A945B3C6138A154175400BE08D0D6DC797AE65B1F7377ABA6A6E0A367A1C07553DFC7F2DD887E14DAE3FA636DAD08003E790DFD0781DAB92F84377F19B863F3D02F03474CEC8C2F5D81850FF1CB0C9264B811978447ECA875030996DE17CF6CAF2334A881B22CCA1F9307ABBEBDDC5621F9AB8C8C785D8570EB9B7701022C20A7A05B4A7694E62B3D0BC3A15A47AA35C9098B42627111F33D5DA5BA9AF09ADF2DE738D03179CC08625E8D33643507E65B2BCB43440AF02618AC114909A3ACCEA4A57F6B3C4AC936AF948A62B2CE671FAC37E392BC0D093BA123CFC01EE3BCA994DA63E67E396F484564F870B3411AEA061BE9BBA2A40539093E5C3F4008A8402A14F1F0C62212AFEFEDF47C70DA27AFEA8A42A9EA5D82CA8484B3220E8AA9064B5FAD14B9F7E6E71D40EB98CD1132F7C9229DBB5D349473DD0A1DDCEDEC0DA9A0611691C6AEEC87535F95E49F98583A7C0FFE948BE7B834609A797DE50866BE97D576153860DCBEAABCA4BBB5483A6BCC03392CAB7BDC104FA4FC7DBF57A0E07B5D5E70FA999BCD83E206784B43D1A11E899146F8C84BEBE3149168B6558B0E025B1AB5C4388381D27711A4275EFC668CC129A7CAB707D4B5F0C04B9A4DF9700ABA4E21A3D7622E33999C232454AF5AA1B36A1D060FCD32A865B55D1179373265019EC3307C51F02E767E9870CCB7BF456D84902B47F6C3A14B7F5690D5D1E5C9EB1E5C9425707B595CF7769C6087532BEBD7F0A8D8E4482358D33317C9FC1EEA75764661F163BAA953305A6422AF50512203E59547B4D6A80DCA3F65BBA42EE6C3F6F3F8A6406515252406C6CB086823CA67B3367A66EEFFDF45CDDBBB5520BF18739FE43AA7E0FF9CD640DFE543C9218D62067EF5A1DDC889B53E1BACCD94A8BE098A55B5F0E295E1D77265FEBD5F399381B027B2B1CE3E977E566052745854F74983B010CDBD2BB973AD75C5277CF6F58B03BDA540E6B37E367396020584BE63ECAB5877F46730FAA2788BB4A48F2B3DE4194DD2417DE2B13979FDA2CD5DA91926C96ED77B90B3099AC339F730FB5F5965ACB8E39B003A31DBA8025B40A98F02572C0916FA386B4676C261CAC365F498E1ED0B6F0E3097A0ABCF8095B132D24A1C9FEA33F3A1DA9A183D4B14B63848FAC0E2233CC0D321DFC664743D93B08A9E90EFDDD81AD615BE873F8D2A84EADA1C541631DBABC1DB65CB9BE534CA984CD52990931DEDCECF08CF1F46456474B881AEA9D166A0AAECE3653714EE9D7FFF3A62A8FA58DE57D02624D571FA24808DEC57392ED16571366C68D8F7D1930073B31373C9E88F5D1359F7C61A06517EC002BC400E0D3D925B758E2EB24857A39D3666CF0132B188EA11FD2515147321ABAF80A56ECBBDB8095C7CF6B14D9CE57A7FED199210BDBEF929B000BF755E5C73213D801D794B5D5C29D25C311E2DECC43866EE1F89E4C3F59B76FD20FC538F1D6E7A1D2890C00272A95EEE5CFCB9AEA4F74981772C90601DC007B1A1C4E3FE3B7688D2290FEA065F5A73E2C82DD63FFBB3462C3F6D39AC9BA4D2BB64899E3F1DF36E77B7C1CFF7C75ECF25083EF7C1AFFBF2596E74C0B02ED0E32C968126666F2894C6FBB39562382F16C53044D1C6E9F23BB86C525F7A370674A54E27F5C32BD2E4FC0D07B93DD006325A73809C5440EA1F9D8332B4E297E45B62C05F4D7F9040C56FB560ACA0F3A7EE942986C95602CEA987AED9C09035AEA4E0D45729B9F190217BA1DC7EAF99A20990D42C8F0FDEB63A75F02F1D84F1BC96A31C0CAA406D0669A3D5528BFA1BA38C122A7FD8C6DCFDAB38CA1839AF1728367EFADBFE10D22110A737B1FDE7AE4A3121A2975D6CCBB08013DE344DA692C799DC4ACD2ECA2ACADE8E819ECAB5B355A5A2B2A924A229F9912852F98F36EE3693EC68FF1738BC5D6793F9DFDC1C0A3457D7BEA73B8B33D548A152FC024F94E1CAB5B62F3E2093C87916FA6E09ECC1304AF4132CC3475D384F031612EA388023DF531498BDCC3DDF4ECBF7112D246CC9367D8118830766495865021923239F624294B148CF09A4C1070D653149B5858B37C2BD146FB7DBA6BEDC637CF427E4BAA528BE6F1FC26E9CFD392A97DA66B16A7822AF3999B1F8D6A96CC32EC2359C30DB1FB932386E6213F1A8AECA3CC8AF6AD67521FB54F583E8A13A4337BBA139A1F2FCC59AB3EEBB19621E4E3BF2EC7A539AC6B77FB22B90F6C863A823E3F093A9CC6E6EF0BA672A64A07686B3E8673E1E793573119159773CA79AF3FDAA0C150195B04E58EE85CA227950A04A281545584E22FA757608637F8DE93A19EE51D6ADA4F30A11BBADB560CAD43C9C0A8C1A76D7475B2E601B713318FFE9189D1565B07E2342ED0536B65E9827D4C8AAC3105A299EAC397BE723AD5CF6F0ED6BC2D023D6227913408C5A570C10D463F489CD27B0927314204D31D34D005398E386A1974B2230E66DCC12D8923280D06191431ECC639C360F96AB616702D4DD8FAAF362C9405661C5D6F7546B9B9A94AF49AF423D4D3E144AB14C4C58668C52611BE6894E6DCE049B7DA76B39EC8B483267309C57713ABAFC185AF09A6C864FB8415DA1A788DAF5EF56DED38C8E363DD47F55FFE388C9B092C0246DC8BA9CAB6838E69C1C9C8943454FFBE34FF33E6DC3EC6948AC0894922172BD7441B8D25FE18500DA31D734E161F9440A12431DBA920968607D8644060B8F033A727175669EF8AD5E03CF0BA1BC42211A3514C296A6D8AD84CA9E1A05924D92E5033310DD8273372531B26397BFCAC00FDD0016A1F12F72D3187BB1CA8A593EB86A868379B3C407FFD8E8DBA764468AF6C1CEC005BBDD91A4E7D3D3831CA8AE90FF7DEF26AE0639439248B55F9E3C1CBF6B0833982D3339AB185F1E3CA3B99EB6539BB6960D7BEC247B26A028E0110524EA8F6055BAA2046CBA9079A38243DFD1EF09FAC4307D625FF6834D6CCD0409E13426B4828BB869226C8330689C474F35E17AEB5E64F43EE8079DB1D85CA4A8238D9D8B60558E44E8A217D8F265AFD4DAB1C014DC8AC9599BC9BDD6581FF034F29F84827C3A8A8F33EE830025C7B7EE1A5D87735A51DC13806D57E76C4035E2C50DA76602148AB750DFA20EC87CEE2A73CFC63C17881692C27DF762FF446084E52DD48AAD8880855D22556C24D7AC171FE3A2CC11EFE6ADB30131110348E5D393E6A8459B171DED361B7FB97B3596F7FEE0639C235E625CB11AF8212FA270A204B281C3B1FD0556C353BED4315FCC59EAB3CF5BE3147A24153DB61E2748A116A737A9EF269E9CCC4BE9088E49E18F2265995CBF430506B424ED1BD84B866CD3CF7BB50608AB48CBBC9D26D8795AD390A654D8C996A179C0B9D691F716937B4D804CA1A92F46261B7B84E1B4445E511E67B2AAE347C6D8339D020BBFF33B22E5843FE4B25BB0E4F31AF46F3D584408B01BBDE7163678B38D54808AA921178F6E4095D7242EAC1F29BC437E1DD0040C8393C1C26F2ACB8FD06F7C066433BC5C196C177F06F45258C882176C680D25A2D9E316C53E0AFC467CDDF02BAA870E38189E4A622257AA07BD3956C496BC44692DB51F13C6D0E76EDC3A4ED5B5DC9B89CED6F532DF22BDAF680E85759E084B8B1FB69BFBC88E800EBDA83B7BC8292B80967B0E2049F981142D935C0BD21C1218966308777DE752B865E7219945D7CD27FCDB6BC150ECF8D4BD729FF54CB5965F4862345A4EF120F6C4791A298D76AC6A5F4D4BAFF245C9B58F886EA2936A307B8EDC3160977A1DC94A887C2F315205DA91F2B14C5948932BACFA1ACA2FFFB56A7C9CB4958BF0C5F60309B3DBD40A6B2A3CC2F770613D70E078783DEFB3A3BF61BE11D60B5BA62798744A3551C2B05FB90D21E600BA0A307CC6958F7E796C9975496BE271DA4A85655F01CB8B75DEEDD0A67F919D00F65489563298459231E344F792F7D85A8FF2244D83D7EF791AFFF246FAF411B1C9A7F94BD48797D94F82E19ED162EFCD85209540D4B5C17949C1FAA8477614F844E35DC1720853ADB4801703D0B30D06CFE616CE890C68E84A20892CC246FD7E4EC4535874CE60B230824B22A504257E7E119E0EB4D641F63162319889D0D3251F512F81C8A96EFE6904A549091BFAB485F07B71CB0D1868562C2FC3BA93308B0FF7F64CF86B6795E43D14808EFA4DCE6D174988F5A9489E2878FDB3AF723FC65AFB0F0EF7FD981949976645164EE121086CB783B0245C5F7875436B333F6519B426507E31E4D624231394A89609FD722F1C61642A375872F561F0730774C146D48CDB33EF536F71D25DC76B886A0D49A94FACC77967B86449A2231B887697BAB1DA877C122BB498E32C4BCE6D0BBFD8FA75E913C4545478D8433D3B1350EDA5C4236BA0CC96AAD20B3D2AB97D7FB45B4D248897157A7E6C422998DD387F5A208733F61E8BA783EDAEFA77A4174DF2F39A2BB29431F881AA9B3CE453333F5660DDC36D95D72AF11832186A11A5E780AF710AFF18C465362676E7BF35B79D418FD17C64A25A8D4360B52300333FEDCD24C5D3E4602B9E5FDBA5B791FB415481EE87110063ED09478C79DB84AFE8A2241C19B035D4315D82802EA1BCCD8AEAE00275667F4B157F943F5022D9E604E239C7A4E169AAD6D27535AC3F74EB5C4A4ACEFE08AE45D3C326A20C53661ACCBB0150DA03CB1A150B9B50D74F3ACFC04187D36ADA5C95127E6533F86A3A63E81314744E4D65DD4DC966F8A2CBC57CB6CF167AA99F77D717CB7D9329BDEDAA0CBF57EF5BC33F5EA2F5517A28CC89CEAE1BD814C7456C9D574EBB9C962F23C047AB36A0B47814DD7D82E5AE217966D75D6AB351F66066F818370017217FC95AAEEEF447D4FFCBEFC9B6C1387527D07923D1621005AA5942742AE83C4B3E1243633E95815A9FD3A31A0F397C9544499D3E8201B19B9FCD4C72349436D1AD639CA2AE5A8DF253F802D5409DE479BD9A99C9A8DB84E8D34EDDC7E44DB7B6E5EFE55BAC03AACFF0E6BA761CB5C7F64A4CB91C2C23BB86803DDC0E3D33991E057D7DF8E32DAA2A79413F828267B240AB4AEC4235ABA52F081998309E08FF93EBB6E61BAFF0524C3710672CFEF951E6F22B2AF10E5A8D441FEE0116A885CBC7FD14E2A9CEDCEF87021DC77D8BF757EB4E402486D62FF9E26A944052933E74EEE8363E7085F51D5AD7FC962280019622F247B7BAE5DD74099E09B009215CBBABF65E6ACE2FBDECF04F4F9C19B4DC9F276CDFC4436DF09C32BCDF60D951FFFC350B9A0BF52BDC7CD8B35904B21399A161E53988B1885E04F278D3EBBA1286EB1AC4F910B48848F719366416E0FDC7251970322DE8515A927164F04DE0A3ACEC85B82E5A8DF9358F6C025DD7147F404A52980BC3F72AFD3D8EF89854C076128CCF60985C0DBCF66F5B88966A37765964DD94EFF2A5DC1728161973417551D3329B2978710A8A7DEE8A8FD1065AC2DB9E1A0AC92D751516B89D4E54353D41D0E68FED78A97F85AA3EDAC0237ABFA1E54F972BDBA484D7A43D44A42A912C0912B70C2CD709A42B0CC4C02BE17F1E0074936F75111CEE71961FD4AF574D1C006746AF3FC49629AAA41570B7E8A18EEC2FAB72B179C4187D81D89E4591BC70753D0DA8BBC9DF9905A9F1AE81895B8E00E374A9864F4137482ABDC0E074DFD7EE0EC89D89360321A19376B4B72EE1DB22547892547EFFC540F4B494BED7A2CC0B783B150D2788D87F015450C80BB90EC70BEBD017E5F63101A97502E009DFD6F3B87953EB98FC45FCDAF79D8DD641E48B5E34793E0EBD348A0BE7DE112AAA0152C1652A3F59B87832E22326FE062FC23F947A119B39ED004A4353DAFEE3886362DD4680D4F9593422B74612E85630B5252C33FC0F758DFC5226E60A61C645D76D8F0C859427989A88D74D507E2637E1AEE80E9E3BFE22807261196975174D9D1983D8B512AFAAB5ABB4288F967BFDFF2AD557D9CD0A71B91A6AFA86FECB84D6C2CBA38CDD078231D8716D0D2CDE50AD31A0F128BC6C552277A4D2076F97449FCEC295721ADC383C75FC558B105A789B15274CF3F594DE4F4F64E24629710EED03EC6770417E0EFFDC902F1316E4164D341FDA56652F06A8BABB67CCEFC213711FFDFC78CE91E25637ED206432F6EFF40CB48BE4BB3FCAFE50DEA77A4E7CBF90640ADF59874481DC345B0FDFEC44FEA753E1B261312D038F7A7D6D5F891EDFD048B1D47F4022F906F340311B7428D1B4D4E721110E7F0EFFEE3ED289432C68903A815ED4FFE849D2B624EDEB234DFD02E490C8A74011BFDE50F5A2B70407C57AA9FF5B16FE5C0B44D116C2A09505E623D0CF20E106EFE3F723F711C23134A3A2BD8E5D60954510FA8E2CD432ED3137C9892824C6895F3BF07753FBBC342E553EBEADAA9BC7ADE8936F3DADE14DB3764941AC56D1DAF2E949279A82EB593120F0651C5CC4550A41DABEEB25B91EC0BE7F78E18DB1A070E68F5A2157DAB8F0F213A699ABA43B28FDDC7DD257B9790A82FF3EF3A0A46838B996BAC1ABB4E3B9F4F15F933142240F676A2A4B537F7CB8C667DCA1330567FA367112F167CF0C7855C16963037962BA15CCA9C7E7250FE71944838DD8B0EC43D10552A6B6833506C4BA0FEBB26B88C7F0AFDECACE6F198DE225C2659199577248CEE6232384B3CC9C53DF5ED7A668B6C823AFFE93CCA75294D09F5B8572F5D47BD53B0C106A6551FDA6A4786D74285DA14C5CDC15739F3533FFF1BA51ECBDB149BDE932B56714E285333FF6230B38B3308C4F44C29E05E54E603E5FCB3EB483F2926DC5561E848A1B93C910EEA397F988F05BE26B3F09ABC073A518703D59E02395AB9DA145A1DBD07136921BE041F0B0D7A173F455E722897C5D63FB21E13DF0ED7B61B807D3498E5B2A213DBC85B618CC835C3A84062F4FBC69CE459D796E5EE794782C66F900DB2FF6F76C070B61683F35FE9101523988B505B3CABF0710BB886FCD311BA4F21C5A18219535F2F1DB12E12DC0DC49AEF9B8EC1BBF551D4CA08B942DE95FA93BA93AE2730FE3EB468A5989EC154C15213E26EC07274189369C0425BEB9714ABF7A5D23CE70570A53EC544910343F07C1C28F48D6D33FE43F5C4B7001EE8517AD3761847ED52441CE477D9E2A308B4A1EF5EEAB6CFED499667CC9C44B18CFE2D1EB0A53F6EFE8A022CCC9A74FA771FF20DBEC02FB91300ADED4DCDE77EAF48CDE5C39AC89EF6815AAB9A4BB244657197C7B3CA77D702B9A495178B56E49CB9B7CEB61A0CFFE6BFF455FBFCE896A6D91FAC883E903C23E34FE157E1FE5BB32A0B2C66896359A238E7629F1B3F4DB06AA8E9C819637A3B574560BB61F8DA87B98DE4419B266896AA63EBA3D62A3E1054112AE596EA8D737D01AF371BFCD22C125059891C4E208335EC9B2D1E773573DC4F631219359EEDF5F946246CFCB9BA3E9659D8B111F806933B8B9CC13D714FBD407B7C94329367C7A1A21CC9EEDDA3EF284ECC0F75F917C2A9DEA78F0847C1B545B2D440214B186732D6AB675DB7C1B086244A9516D75A746D93309ED92EC262E4AA577A38848FCDDE72F380E3E2EE617E0AC08CB94861A0A80C245E2CB07F48A0C06B0DF145C511DB4109F739FDF969FB5C0FE347FB1ABDE3D705AF6CDE3DF44EEB4326D3D7497AE2ADED7AED4EBF18ABC0B7B338FD01CFFB32807E07EC759E4F180086E12A6F7E6E6CD92C2FDF4F743D81FF3D65C266095D05800EBDDDEC6F3319EDD339E90035DA7F1D51461D6FBCD4F3AC5D66A0D85AA4B857DF6AD16A0289F5E060D3F52E496D88111FBCBF7D4600F22D19602EC4D45F95B2870915BF50937A8FA59BAA9073C34FB696BB364B1665A2B5DE9D414371A64CB15709F3D0CEBEE5501DCB5900E39BF46A1911F1E504F825FD7211E273CD4DD8C451D48A08F7B72C50C6B999BE776C18756E1DF41ED96A8F2199B2EF2589A7FBD4154BD571E054A0ACEC1780B182BA0B398BF4DBC0C21BBDFBA2636272D1863CAC01D24C5B8EF12CC482EF641DEE9B11D32215B1AC10F92F07CFA5AB1B1E95ECF2E54FFCFC7D6A35C497478EBF07E54817CF44951A8FE54F3CA35A5C8F3F98BDB68E540951BECA05B6EF9D8ACC531FFBB30E366BB330B613DEB9A953AB28E5447E094CB7302E9F01B374B498B9143DD87AEFB1431CBD2B2169E7803E6D63779FD69D570AFA11F76E03E5DB951310A5212BF46E9D14814E8D2D140111E371C5FB9843204D4C51CA986593C1B9ED65377F678277B83AB9FE5F2964A233C4D3449532B2C0B6B605CDE09196093D5FDE5FAD0D0857C970C542E99F435929B77CE56AAF17E4EC4D70840AD21DF7883EA264DB1B74AA919640CD6F486D53EFABAAE99C0BD0978F20C6C7F230695C412845DB828D5A12197677EA375AE00DBAD37A55B851923F30A878E04397336C4110C5D422A4B6F091880F61A58C9FC78427B6412410F6743B7AD9C1B4A37600693B995EAAEF3EEB264C2DE1493CD1ACA64FB9CF5D1515CD4D2EFC91ECD958EDECF994E0EAC37A9247F409B5DF1807A1074B54CC4B3661062CABFBB1843218667E5F7EABAA9690F0895C23300ECFA684032245B991C6B0B292439A1E6FB682D07AEC4F4263708EC7DF823E0838B15FD22EAE768D0BC23773880614AC9696A1F37F048476AF79E725BF206813BA6EB149DC93D395E6D192DFFE52EED229D17B2AD19F6B7464735AD16025E40096D00FF87BFEBFB5810F1E61570D960B8E9FD583DE4B80ECF666B578CD68CF5DCD2FD2C01399E3A9DE0DB1917DDE37BBBB919ACE61F93E2413E6AE8C9B0C44F10606BDA347DF064437CD33FAD5F66E7958B98F4118929D9CC06B6B5262F884B44EADBDFC0C1C79680D63403F13E007B2A9C0BBF00356A8C565D77BFC657F84AF33135640246069FB599F442740F13C983996857A2D6A389F7CEAE4355E0B6D1A56A5804C71BB87C749432832EAFB86D473D9B269E3388A09D8BBC6596A61000E5809860C4707CB3E359371A12E0A4921DF1E33C44665DD17FB739BF22C191D10126A05184C3A39F638C9F40F4975BD7EFB92BA44D53FCE48C1230E4E89C96A780E290A501FCC51A6380B8CB07A7DCAC93348EFF2175FEECEE359B090258628C28E90B9713474FF32C0ECA86FE6102C9AB054945E934F94B699B5471990BA07A217EC5DBFA258BB4FC685048153833BE625466340F9F8E50F2A6D3D0DCA56A1154FC85452AAD12568C2E92DA6BA52E81B9FD8A70C4194404CD71A9436A2097AFC5311C486F3A1B4F17A698C8C4A1084677BF12C104C9E26462DF7EC0EBBD56F5F642CE22E9CCF0F0B0D0F8EDDC4E755DB64D39973680364CAE4A05F149DDA0C41F63880346F04D4D00F92F6A3460383FCE05ADDC1E1C79EBE5E267B3BA0EE5A0A224477EA315CBF73C9BCC460FD9D0CA3931A15F193F9084D2EE17EEE07A7203B85119B034F28357A53EF39A61BFC7F3A4263EDB5E5300CE34EF57603D215EE90B8901A51BA0B57447A39C72C3D5454442B0CBDCB2519D6FBB63E93EA9AAA3F33656D2911D918FC73F6AC03AEE1C9E8098203C4CEAB86D34DCC2EC5E74E056585ECFDBA978090089892EAE7DA5165BF7CBACED561BA3FAE0F92F544EF6B3C00CB508A37CE2B1C062E198A12253B75AE6EEA1380DEB4C3A11C926558EE38C5ACBC46BE1C0F18EB351CFB693351192BCFD64FD24F4E10D697F22C37E4653B7C98350CD81B7AF2A35C44969123F7704288E0D39802292F2DBC7304AF2B401FCC29549001B0DC4E02D3A727629F0193DF00FCF30C6198D1A9B89959CFEE80A2D4163429215198439B2746F44D52AAE9A32FC154FDEE4CBC8C5D5320EA92A3E886C34C44B59B1365CD3C75EF976F0FBED85DA439565E02470A87C2491CA9CB713A60644095D516C1BF1D94D8AD039DF6E3A226A08CA1EEAC7EA4B1C0CE61419B8BB3DCDE636317730468BC4F01E5D7F2AEEA99995D30B57FC21A613695FB09A44A91A109017A4D09E8E04CCF523EF49B6BE36319BE2020C00AAA5A19B3604A86573585FE13CAD8B5CF5DF48EC3284044874697F6407B5D3D24E092FAE370AE9090B80033CFA6A67915988FFBFCB5DC698F586F62C7AA647F3A29568393C49FEF935A062FC531F0838366DEEF24444F7DEA1FD9830A5B2D8B18DCA56026BC6B45D985131D7FE9D4AFA945CFF5F621EE20C0D319173560144F2BF363DC7490E86854ABCB6CD5AC8957163C29E81D8A1F58F44EA8E1CE41C333C6E73FD628B5CD891D2D3A4261F40C5C8EF58C6691BF9EA5CF841082AF61E094DD5827132763522B9597F54E37EECB895DF428B03818736EEBC768712DAA2256E17C9262C462C173FB2607560D07778FE264DD43946BE5A9A9CF34E3547C17F383CB88B0E6945E3D929B86F79A6A8951A723BFD0D1C6074622087A4DBD3BA7BC2961917BC501847453D653AD8D70FA817CA3B2ADDFCBD3DC403530560037D412C78B3211075AEEAD41D8624286B4A9A154490756DC36A5FF5A67040347FC2340692BBA0CDACDAD142C1DCEE4A7E67C47B7CBF790A19125CD8E40B352E87399F6FF3C2F31C5588980FD867E7CBD876EA975C48F41263335D0BAB8803B4B06327471B8A2C582D0E1B665D3C041FF5368D0108E15FA7B58F0779726700F95E1B1AFE7FC2284B310FDC016D7835033E9C0FDB720FB82C29499A069E385B41361B3077016983DE0774825009DF8D7B2CD74E65D29FCC031FD432D29344B63255F508C4CAABAC52BA38C8B04719797894584F7B675A245734FE2481A9FB271B878F8D2FBB358052F2A00A6C176D483B1CB2A6B0B6D90B37AD02679A236AE0D968E6604E81A181CFA1CA4F7D8F7B8964C8DE0B62457AF507BAD5425E2116293247AD5037E3949310FC4874797486DF596DD56131A8CB95814688D23200610DF2858596D2D2615E0D92EC8A8651EDE5025577196F95454C79DA7D314C1B7FE52440E64C6CAB8F6AE370A8EFE0E7B4E9AC2F47E4B22CA8F3A05A7C30E8E4ED9ED2B0C6D83FC8EDB7B8EB85D959B12906C39D45ECAC8FB5E6DABB0ED4A98CB330CDE0114C0FC46EA85E442885F6908023997C779709A777A7DF207A9263C3646054D066FC81723C42C014351B258CFBD50E49DA4D9160556E78B79FFDFD71BA0E35D94F2C62C53F1FE3B8AE48953EEB51FD435D2747EFB263490932DF7D67B383857919744A0030D1D6C2D7E4705AFFD6C7BA1BA9A7121485B66EA70DF86BB12B4AA57B1F5F54740018DE3CBC93BF4A26D16CB1701B464E08844D1271BC796F50A02A8FEB104D89F42BCD852FF490170ABBA550184E3F5792CBF7E9CD1FC587608A24AF1A67455959D54C92269F8CAAC5A0943A1DBF1D4071B4BEAE1E53CFB51A796577042D475BFC9AD584A850FDD0CEEC671DC8A230F84B590C257297468FA0809357C6C0B001E322E4A06068BFAC945470270E0B08AE75B932FAE9E61281AB1C6CFB4825C868599AF3D91CE2653571FFA0C3EF5E744F23033C0E29D422FA4088447325888AF012863F9EE59490BB4268A393D82FB9CBE9A25A4ACFC24591285C657C1DAD92FBB123719371A185FB6B1B2E9FCDDD2C0B03E4048B6719F8DE338AEC69864A5CEB06C5582A6CE8775DE398F1438B6D6DC2B0029BAA06CA1FDF7F1A0321F8B30E343BC95CA545A3E6F123849CF61BC1D29F5BEB0BAC5BAFE0B5F27B505157EACB9E579B2901F28CD716447DC5E678D4D9F25B34FBF1530529EFBCD678C88D24928A595B7ED87A83880AF2BD9A3B2C23019DC0BD50ED6CFF56493E0E8D28A5E8265C1B1855CE08B1C4F14D0CFC03C0B9FD65A3A6A1F35649A8F6437EC8C5E6E58CC949232CC0CFA023829A82715A8D9626B1CFCC31BE1ED49036CA89C1AB70009206047CCA322A5349C8B352B3CA96FAE1D869E43AF0B77377C8E5564488F78D47B4999218DACFB86C0C3F330F6D33AB89B6BD0B7052BB19916F8AC962A1BFC05E5B808534B6FFA02E356B0275D76496BB039503AE414F9FC947001DCF82F820E8EED66B8DE43EC273F2972DA346CAD2D8C15597D710CA5781E9F81EFFA97E062EF95AAC1EAFF7B6A1ABB35F1E8C6CA34F275766AFC7ED7AE5D9103319EA60B366FAFC2AEC687A4879C656603D0AA8273F8F7D86FC9DB184D18B0D599D0EB25C6DBD2FE9EF9EB0E4EFDC4BB063A6C5CFE3F4B6BC02527BAACFF3CD7458DB31CE7FA17DB5C011BC4C1A2BED7775C80F9EC1F5703C94C8FDAE6409C7A1115B7E8EEC8799E27A33774F19315766D3307E445266F3BCB94FD95F7D9621E2975C83EB40082465F6796B04FB7B16FC108E7AB648F4BAE4FE00119396A24905C381B53DF4029B97BA62B7BA7FBC288B65967E77D0CC914A675194F6FCCCEC77BB0488C65C88606C924D66E73FEA8E58A90B8E506F742520B14316497338AC4BB047BAD1FB6E746BC77C49E16A94F1BA96502A0B3FE1A7CA3E5D3079471353FE394E2FC988556A6C81C7B5CB01FE03223A4DD4F1A360B25C9D62793DE7AEE19E9B409BD6B92727DC8350BB2E427DB73A6C34B1121A8AA54AE1FAD26DD1EF5DDED4B89F009F2AEEF98F8DA7726940B3BF1786994E57E589EC3217DC37A756926CB6B0397D4CA9CCED49699FB7912167330CB989C8FAA79AD724C8A49390315360228E5845F5AE3E258F0B9E51849883EA1985A36D8F32B12519FDFBEEE109126B05EDB21D518E4601A6DB378E23AFEE9B528F38209EEFD8F78D6C547CADAC0F50E15C5B5191E93352F3D2D1312E9BF0E43A4DD0A8024E593741C20646A511069BAAC3741A442877F09AE0A65B99100DE8C3D9E1B4F72D7C9AC18E3A7D512BDDDE05EAF58AE939206AB606CCD60794347676288D3528642E9336BED7F1C6BBF6C42C267E2B8A3EB87D5F7E80789A5A3FF35FD1D687F8DD91723C23EB51AC6017DE6B87B4A1293894E988D28564007EE8F8BF931ACB411B2DD9705D502441CF7B20BCCF399290D0DB4C52E48AEB8002E394701B7EE448CFEF76A89612D0AD664D8DEEA63F011F12C19E53AD287E388B7161FBBCBC3B6958AB56C7F5AEC4FEACD4C95571D78F64C65A6EB2EA03A1F47168369B19FEA78B7589604C4DA76BF2C9138A8798C2369C0FBC908BBC32DDA45BFDAEAA815BB9C6F7286BFF6AAEDD4950B6FC20F6E38A57B4CDE4350CF9D6F43221BC5D0CBA23EE80447437A0AE2680DE548F42E2B602B4DA588E94F121C305CEA145D081FC7E6D022CE617A1ED9EF709C38626A1697EAEFEC41EFD457A66C12B681300BDCDAB018443B0B452404D7697EEB9CD5D280654C17E7292E70AC029E7809649EC85F0685FA87329DBB28704C250D231273043950A331F89004005D126E27E48B57D91E701C7090870D2672EC2B79BD07B0AC5D1795214BD78979215F15AE19B354B7259580AEE76DEBC1A13D181846296E27A5B0D73805F85D66C1A60A461BF1F84D5D70FB994F11C393DB409FBA6F9749A12B6E42ED4BF8A0DE082B716D9BC4ECB0CBCA139E006295ECF96BF5BB068E994F98EB231F7233B02E43C52C079C7BF2EF3385515D508BBD370CA3B147FE2DEE633440045566E2354C0B99955073D07F1FE8B86D6E92EE222A13F6BF830C90987A58CA71A006EC54B6C0B388FFD447F2148F8FB61843447542E66CB72F6CA38C083FC63123BD7286F8C47FDA44C1B9C8D594EDA1887A49010D7C6A944FCEFA8D51CF258BC2C6A8F694BBEE42FD85EF0AD75B10349AED18A693846BE220EAF48424291E41EA0DB2D56F9FB345F81E9EFCA12AD5B03836A45F860EB08C9FC287AF3062FDB5B1BEFF982173BF578FF227A2D39E997AB8ADFB4AD52DA687C6D2025C86D755A494FF272FD1820A632D80BC41FF789AE5B2A0297919E9DD3688FFDC85CB6C912A209F83470404EB0BC1DF052C41A4D955FF0557CCE1283FD606EEA4CAB654585350E33ABE0AE982EB85128CB5E4F2322C89DCA5046923B4DC87F8933111C0B9A952D4B2782CFF96D3FBEF18685006BBEAEF20F6457E33B12C6D4ED1DCD87605689DF92788E979EFC5AEBE2FB3A2198EA03C35972CA4A908F5F2B33247615D82C7E580302946FF64D3D6EDCF62524FD5B75B7F37CC99AC1ADDFC3EF82073CBD1CDAA486B3A24B45D7BA31C57C4A26301FC8793989E220F915ECD484FC2AC3B2AA88E4A55900BC0A3640019094F9299B613610AE27682C8CD9B8EB391DA908ECC43BBCB6CC1A8B14B2C196E3B09FC27E6AB3B47A9771D24F5B9FE35E8751F46F04BCAC2FC837EAC5679B440BFDF1579DA031E5629F9C87EBC3EFF6BF6C999028701E9ADB244753B50D08F729C064B9370465B115E59017641938371B5B54A622A64A63C7F91F331A9969FE095974F759CC03BE2734782B745159BB6F85934F9114809C9CE478312B9A1CEC0CCAD95BF792D6313406E6A42BAAE7B4ECB286F75B3C5AF9B7A19CD77483DE289C46FF28C9DD253F7D4C8FF51C1C93EA938DF87D71BE35F99C16816A05291621C697B267F5F5F00E7693B8A0F9A3F673F6A8CA7A8406AE04B75A16948B37646208DA9E02A093EAFDFAC62515D702DF06553677D2E60D0E89D50CB979D963A776E7C9DF08A782913510D63853E40B9FA88BF3D53A68447E505817BBC46F9D8AC2D70C614CCA346F447D116066EAE395F28286D0D5AF7FDAB3B69ECD69B88DC9ED8D3BF668403B8FE8F59F98338E1B18DE21E3212908C2E12D22FE0B948E41B999DB3B2588F088C3AC4F678861ED6EF54C103A8CD33F50B507D8DE8A2E49C239372ABFA1E24FE9081CB2F35B9CE9FB7BF164D33EEE314C4237E6B8B5E2DBD954450E81ACB67CB6E0DCEFCF69DDBF4C04CDBFF4E1CD01DC22498624841C157977013A88863D9F04CA1424F19F54AF8A2EAF499B09265581D0356160378C4B2F0BC08A18404382960027B4A9B9A340E8A1F8F480D1DB6CEC10F4275F52D7618BF97C0EC632296F464CDBD875A8BCE6F49D3E88863AB1E4CA9FFE0574B6A45031624D60674982D05A2C458365F0E9B3880CB76BCCBA7EAFD197AE814AF4CCE7B0B48CB28DC5771665A4DE13E03EE78659883D11273669AAA2612E165F03FEA1E41B5B4E543AF264564EA28D21286014AAA4531C9484834BC11E0BC223047CF6C0F643EBDDAEB220B92FD1B7251B58269AD6F15D608718863465D5AA98FA3AD7007A0AE555E82CC4EEE8C26DC8509887FB6B87DBFA40F8EA3ECBCB7224348EEE27E0A3160BB001FBF042B32A2586E1C3401651EF4DAEA1D2C2F14A3D2419FD31EF581244A597BA08955483468B1037EA3B27FFC5F9F6846433710831CE0FB3F82C5BD4BDA0FDF769387298C529EC23F0E8F229B0E272CC26DD5681E8ADD453E5060E76B484043788469DD19CDADE1D8369FE914FF6EDF01280186E32DDF7C6406259243254D2E5FAD02113AE5F7978960AE59B894E0EF58EC4C01F3FEAD19421D2065285DE72E9DA7569654B54E2CA1365AEC9D2CBD8789B40FBA14F312CD65900044C5BA0CD55457827DFDC9BB14FF21FD2B9B40DB1417DC32F32F1238833C9F831DD3FA6468670C8CA805DC855DDFBFD134D233D82744F5A3D6DB86656FE617A52EB7848423746D77BA18175D3819C11717003C58CA6CD9C3397CD94C58040A456643468D961D95C283995833645C00EC0BB4C37B8B060B71C3644BE42A6A7C514E110E38FC081FF3C53A578EE79EAEFDAF6C4035360DF7C96984B8829D646F5C3EFEE9A6CC7A4EC103D07A4576C0F2C849EBC1403502D5511B122A3CF71FD066637B9508BB34FBF726AE0D092E16FF0AC4B8B580F312EE77251C8143D32BD91AE32822D7E189C98FF392349709836D5BA65BF7AFE2F5E9FD3EFA6687E51D718E6D5F75EF8A12F1792D51023D7F6C12FE66B1D3F0F753C671149F9583CF7C77330A02516E297D15246DC2848FB7E6FB1CA0B6BBA2C8F1DF3E3A0C309207B23457D528CD27648FEAF61437DF42C0477452C310E0168C256B3F9E5F1F8173AC1DC1DD7D02B4F748935EC829EB8FE6C8C321B9CC3BDEF75464E00A3BFE61F07EE0B3D11DC22A064D4548B00CDB9F5CC6E327AAD2AAEF9146F6AF4486B39B0162F1C010785E537E35F7A903BAF7CACB8F8A568087AC23014218335B48846917D0C94D2BB509C326B79EE9949E72DDE40688BCD31E621ABE8FDED1C1542CBEB12C275DF9351CCFA75A5FA277A01DFBC15E8CFE6F0E0FCE6BDE87E4F15F21B8F0BD587BBDCB0F5A125E177EBD453CE3D5A96F5EABC89A9ADEDCCA7E5DD55771ECBD6563A829EBBCA0C4CD594B5F291A1FB7D60DB64696679CF40659515E00FA7F966513A77B3567C10D01ED2EED8535AFA03E7A537FE8C8056F55F55F7FA00F0DD30029A3DD0A9752851DDBA345FBA88F0F4246D06564EE62D9CAF6E9D4D5D8E511143A6FDDF199B0537FC02E6A1127DAF5E87944AA9A67BEB8D51D3E2D16E62B11F46463E187DD26819A2B67E987BD3648F83A6B57F4E4A7F7941BBC6F668050D87CD19888A5DAB4B8A343DFF9F66B6E96A4DC3B4E7A062350168AC325B3627CECEF47AE6898B6B31A3960786FC389504C65BE071B0FC4293E292013D80274F45E4FF266B171F744FE6A1627446DE60BAA0548B3C181A24A49D634932DA947BF4E02535C66EF5451285740DC8AC78D6E05262D9D01DCFFF708B53042330A843B1BF674639B1FE39AE7D3E22DF86F45266BAA99B6DD07B98130DC95946672AC52D5D65F6EBBEBA7AF33870B324D0B7EDB4AD1F5D088A4B7E04BF1FC7A23912876CF34181601FD677182B41E6C2DB29A275AACF990ADE9B75D5CB00B203F48CAE438CC6EE8C604AD0941CCC1452F36D9FBA3CC0BB50D8AF0211A8AB3B2186EEFFB81F2C26EAC7DC0D060E48788D00C79DC6EB89A2F045590713B3A044C2D0907F79076DAFCCE658C82A5902F537B0613ED665A82B9CDE61B657CD0377C4100C9291C5B2C39EAB0E779A80481B93CBE97E49DC1E37566BB4A9ED27BCCB0564B99A19BE43DA8FACDE807CF92A804C32417462480E43090719D0036C5A0B25CDB37E5427AFBFCBBD25E3C5F95A2C95D21CE6F74F0F4577CA0A863B4293EACE96A46748A8D80CED666ADC1B0DF3732FE44026DE8116E6376B82F1E27FEC2865793D05C84475070F4FDB13F6BCF12BA986E60CE82099345820E70AD3A8C38DE7F8BD6684EB117FE507E35E6A24B75A9EEC422000E5314915F7CC034FD93C8D90AD4C76D5DD5E3199A858564DD9BB7ED9384F6E707BED1961A43E2CED90D3B5C852A09FE6A148481EC305E78252265B17EFB42B5F4D75973E5EF404EBEE25754E7BDAEB15F7BC883E2B26C385667906F0D97D1262E7F00FF9A73B3B35863494775963DCA6DFA987C2962F3566755A02E886D3B40A9177EDDA685D1ED71DFB0FE1B4223FCF558FE4B768C0DBDC8BD8BBD02ECE3B4A2828AE99E4E55D02C830A53142026466FD46BBEE8C1EABCA589A8B124B661BA7D53C23172DE9C6F6F47D639DD53B019BD3813EDEB8D8F2AE6CECBF054B1DFF94AE37B6CDDF052A305A5834273CEDD692081D61229A9DD20EC3C73B19A194D65D504DB20B43374A57BFE59949531B8A2EF715D972DE8501F35DE969907572C9C914A52AC2D763FC8301F2D527C042A06F5D3F8FC42DC29413CBBA198DDA30CBF139544F090AB92B25FE81075B478CFA970D4A67AD8F20FE53962EFA05F5ED2EA6E154CA3689E7DF30F082602EDE4C3DB7DC1E8B5D01A491F53F9C9AE666118277108D65B73482E451F693B67BF31A10224BCCF7E3778DBF7CA45AD3E54273F236DACA32003C38E46E24EA02E4B67998BC2D5C221094B9B311F650DDB14DE78B2B10B3EADDC7FD770E4CBAE43DB8BB2D31FAFB998BAEDC87BA67FE1F6157066A6770D32CE322E45FF21CBC5A4C37040472F006CD80C807BB2223A6C88597087CD6CD2FD15174962EC5A56C4AFD053325B48CEA6D73BC15B1DB536A6FE14156F404D893DC6C06A880334FD613D15621054424BEBA935AD3A40D71E13CEAC70B117D04F4930E2B533269F70DF9499F99D280C422C9B71BB1A700E67F6F6106FCE55F3C14793FD703A9CDC3416D5731629E484F48576695B2E4A8B06AC6028D993EF547E2969F3166A5BE73C24D334FF96A3DC054B8CEEE4C2FD6687C803FD899C137F423B4C7395D29295B63D62F4092B7C9B3E636C6D90775E529D5FC678B367FFBBC05E9E504112756F4565EFBA337C129364E6E56860769D71CA8C52250DB54CA4A541CDC006F903CEFD6DB1446FFD1329FB54AB04FA75CDA29DA1189A74B6DC10FDF96D66686E68DAFE8B5CE791EC68716C921B15681F40D20BF83023B9EEE1C5C5BE2300D5D07F5B786F5F43711D4DC243F745E41FF90F8C78EF28BF2B0456D120F9DEAEBE3DA766ADA395A8DDBFCE25370A6F25715D0C1C1CFD8926208CFB023B02F5A4A4213145A8895D25E9C96CF0B325024194F49E0B1781DD21CEBC53484F2A1984E03F640B591F25BB2CB67E4C2849C4EE4D05D8BE5D8FAE86E71E932460AA43D20BA4FB9F3E202F3EAE7C9353AB1F487069B5A0F769D3121EFB33E43CF37B6492467A8522A359653D6B3593E2149FADB1849D08D13D7E102E7ECA1F7C925100423C1E18E6E4CB78C9319AD77BA16A5C729B700533DDF7AA7779E8DD761766DF5734B4FA922C1A0C2068379E1B6A02FBAF373EC041EDD0B204287C008BC98479249DDA1BB38CEB496C9F15F2994EDBE139928F8648F56F168709C0D21637BC45EF7C39236A56CDE27E7EAA7D6651586D5C23A77258CA4690C4A9383A8BF27BE81E570FB86D53A9E1CA52814145EED557DEC36D6DF09F3B3C14762F6D61013D41FB6063846CC5119A850AF950D6BE9AFF504FA8B22873B43829A97F380C209CDF7BE48F579AD016658391DAF4CD02821C0B31E5B9DD60D446EAD43F23A1FB28DCE53D93CDED73735F143FAC5C84758D713F7924E92D77B4BCD49A9934AC218D460DEDA28EE25A497CD01D7570781D2D9789D5EF03C89F4890F1F6F6DF9846140CBBD90CC7524F13FD58BDE6C2A6968AFFF969213053A6166E1ADC0660268DC6D12C223A006877E9AAB00C44621F1A319D058A7885FB0821816124B6F8FF0D6097F598F1DCE982D7072B4F04BB8ACF0C74EC1EA5DC1B6082356DF3F84C3A6B640AC288F378200DA1EEEAC0E0530F3547A4016B18AD754405E9757E2CCABF8D3D883BA0F8818AA3867A07C8D88EE9A436A65CF8F505DF039B917F8D797585432908F72B06F3C893C4C71C62CA42F17027F01B9EB4CAECA4B236ABA5177B1AD2CE2835C3E1FBE5F037CB4DE3D3EDD64AD8060AEEB6238F1E241F9C790EEAAF33A482C5687BCD7D83ABF02DEC875E41AE9FECC15968A36460CEB710E4A99684EDEAD153BE33136BCDBCFFA20CB7C9931352F46F416816BF5E5BCCE89E827E852E428CD31BF5D99E5698B53E70CC65258E438CECA4B25B81E68D3099AEEFE9F336AC3298248566C394C5C194123FA07B8FED0A6A5CC424A888681935B71925D0E87B35847F73FA951FE2F4CC57E20A426A9C5552AABA0ADD3572D1F1242F143BB03DA881A362F54D4CC46A9CFDD9BF5473DBB51B444666EF4AFD9DC6FBC63BDCD8C204DF0FAA2C6873DFC00F62F64B1FF34BD58D34C5680F653DA458A8C7A9441009A770B7323A9FEBC984EF21997AED362C8D255D28B0AB2A8EF643C17C177D0FF6A4B9A5D368E0A3251704709526B2961843514B72D99163BE01FBFD48257C10909D0B93B2ECE5CBA2519CBD46863D40152DD95B8C8DB104FB8CD8EF52ED39F02AE8EEA93D284F8C7E6F314D7D9706B55862333ABDF6D1638B42743E1563E922B3A2FDD33CCAB68619F2C812C9288A8911CB3400406AC79CDAD52ACD00B28EA05771F146058A890E2D6A9F173F2A945C752CC4A64C8DE9AEDB31262EF64457B07C536521609BC4174B47186CA26238C3CA925F3551090BC2B22510D8A66253010C00F76A2C871FD111F6D3EBE5AB7DD8B71B1905383E13F5CCB718F3B4E7CB6837F50B656D4A5FA99282A088209EA708D4CA48A3C43D02D0DC79B344C55206A8037F686AFB36FB7719CF35C97E8A6B0E54FA66D1ACDA246AC2ABF0F225A6C4E8114E786563B5D89FBCB2F440F509A0120D8061FEC0E6A376A992076EB34B028573D4EE3E8D2B84BBBAD6C772285B2318D066702358E2F5F0DA0B7ADF2B7AE04C1D3D92750D007C6B21F2065C7DE80F492517E39437BAB90D8E9210328229FA648AA847871C62AEC37A09A2FC03F7B13D5C5923ECD144666AF53492E31C9F50DC5FAEF55C41AB671821BEF0F8B4ED0E9DB766E28502B50A991930B689F83274D99C465E85616E931B5DC0596E814BFBF8769FA455BA466B3A54665E72FE0A1B3A8696E1D6A27892AEEEE372AD43DA6C9DF95D2578FE834B3D2F35E9E5A211E17EC97193E9FB8EDC28AF863DE7EDC31ACB5C80E1106CB481CCB5FC09B17714AABEDA5669AE60478FD5E421BCF056BD0B56BBEE714BEA394808458B68A63C5C233B1F7A550F41DE420EAC4D69406C8697E4B1D9003703110C920E6BA2A09A95BD6BE87C3BD3783870FB9440283638DCDB462534EE6FC2A3FF0FAB7EE65A22306759F82FD7C7231425E16830A641AA7B4AC11C6A73E269CE6DFA0EB4C40FCA5038025D40C0B0005043437B1912102DA46B4169FAF61CF4A10AD996A3056BE6E6E3677A285C6768E3B3D93B1530D7F476AD5774444A004A5F1F1BC90B8E58B3C1170FA767872E0680EE1E9ED3DD9D3ED0CEFB52F31D893E8165D5AF10C311B496879E619C4818B7217BBCD8F2E19211F934BAA4610D5658E563A1CEA40E640A48B0543ADE5434E4A8AEB504632988324DBFFE2EEDF8A045BF387C682D21144B6C63B3CC61DE64FCB0A83AD551781F184E544C1DA8F4534C386F59F2F1281A112A65446203C7078997BA2DAFA1C60D1B8AC072C4712E8D24B70AB3E5AC15A535A18222BB3D8575063D058BFCA03A64C77A9F33D2CBCFA89B4482A915220177310D32496BA1F551BD322FF274A31FA03EE6762FEBDB6B9BD6DAFE2A09AEA5B5E206E82A26EE254A9EBC9578B00818993C7B450A0313952138D5FF51634497AD21272687C4CE447F0B6700EFA052D6993B289E01C5E96ABBE48831032C67665E89EAF18AE34D59087A87B01F838F98BE4DFB377AF4F81AA1CFDA41C976178E2F38AF8208A2461BD4892FB018B7DD979BD8176B9BC65010347AAEBEAFCCDEB89BE'
	// reason := 'valid signature and message - signature should verify successfully'

	skb := hex.decode(sk)!
	pkb := hex.decode(pk)!
	addrnd := hex.decode(additionalrandomness)!
	msg := hex.decode(message)!
	sig := hex.decode(signature)!

	ctx := new_context_from_name(parameterset)!
	pkey := new_pubkey(ctx, pkb)!

	slh_sig := parse_slhsignature(ctx, sig)!
	// slh_verify_internal(msg []u8, sig &SLHSignature, pk &PubKey) !bool
	result := slh_verify_internal(msg, slh_sig, pkey)!

	assert result == testpassed

	// Test with PubKey.verify API
	opt := Options{
		msg_encoding: MsgEncoding.noencode
		testing:      true
	}
	cx := []u8{}
	// verify(msg []u8, sig []u8, cx []u8, opt Options) !bool
	result2 := pkey.verify(msg, sig, cx, opt)!
	assert result2 == testpassed
}
