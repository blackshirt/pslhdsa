// Copyright © 2024 blackshirt.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
//
// Test file for fors functionality
// The test material was adapted from the golang version of slh_dsa module
module pslhdsa

import encoding.hex

// Test 1
struct ForsSKGenTest {
	skseed      string
	pkseed      string
	expected_sk string
	idx         u32
}

fn test_fors_skgen() ! {
	tests := [
		ForsSKGenTest{'00000000000000000000000000000000', 'ffffffffffffffffffffffffffffffff', '5119e92f1e3a5f02e86b2d2fad9f8f12', 1},
		ForsSKGenTest{'ffffffffffffffffffffffffffffffff', '00000000000000000000000000000000', 'f594fbd328494c749789eefe1bf6674b', 1},
		ForsSKGenTest{'00000000000000000000000000000000', 'ffffffffffffffffffffffffffffffff', 'daf49383606b6585fcf94a0d59fb281b', 0xC0FFEE},
		ForsSKGenTest{'ffffffffffffffffffffffffffffffff', '00000000000000000000000000000000', '6dfd40cea244d8aff8edb9e252871c36', 0xC0FFEE},
	]
	c := new_context(.shake_128f)
	for item in tests {
		skseed := hex.decode(item.skseed)!
		pkseed := hex.decode(item.pkseed)!
		expected_sk := hex.decode(item.expected_sk)!
		addr := new_address()
		// fors_skgen(c &Context, skseed []u8, pkseed []u8, addr Address, idx u32) ![]u8
		node := fors_skgen(c, skseed, pkseed, addr, item.idx)!
		assert expected_sk == node
	}
}

// Test 2
struct ForsSignVerifyTest {
	md            string
	skseed        string
	pkseed        string
	expected_sign string
	expected_pk   string
}

fn test_fors_sign_verify() ! {
	tests := [
		ForsSignVerifyTest{'9f86d081884c7d659a2feaa0c55ad015a3bf4f1b2b0b822cd1', '00000000000000000000000000000000', 'ffffffffffffffffffffffffffffffff', 'dfb10edf76c996d39e0a64ea547e6bf37be32231fb8fa5855787b59feb19f68edd43b77dda873d87be343a3e8488adf7f11f7abb4c3b7d876c199af0e1f9609bd0f9921906435bc756e2f45c52d71d9cbd4c471b8890a23de73793b80f03703ea86f61e178dff376428abdaeabe7de1e158953da03252c7358fda0505530ae974582ce42b87286aa659946dea36497194d5b3f30bc9bb03ad0df6704984742a8d7b29dedc1c74bc93d444ff127a5654b5dbac0497916f774afb9af58521bc67e911a0fcf5e2be5f12a753d387d3b9f97fddff3cb2eab81c4e30b352d1490328bafdea2acbe271c89625243ffde3e9f27eb8d44782384d804568ec8f0a22be5c3df9d79e0f6c567550df5bebf2c15982c7e541ca04641145860e762525ba1b7f2290e3b8a8a1c2389863a8bcc3f1cc800791abd662a4ccc51cdfaca3df404164391f13f5934b8133ccbac321515f316d8d95a41424ee42fbb09f08a8850446e3a4a0f1224831b8679001a630cf9242b49b5a83e6450612ae2297ba146ff38f06e203f6aa2e5fa5941ec8e84720570042abfb486058c75138e2156f22926faa1a94693ae3472eb4b3b5f87d1109c528a0e5f3ff021c46eb97b7e2e52808192f1fca86603d48b84ef0b92f7a712b853b9030e5b83574a4e8944329efd157381c6dc2254140c0c2631d74538d8fbf76d8bb93445cdc3ebe9c73da78146afb357b2eeecd78b042329ba911c50ccd4376520d9687b4cce878961cc049c29e251a9b90efc63e2e27e918a146679edea2c73d6d38cc8c5ccf2ce715653490ff5b986feb93afec5ccd8c0bbf21a2d39b94b79fd1615466ca52e19df43bd67d634dd962e64b704996b9dd892959f9707e872a352fc2d8e17a143780724425ffd4d3288a8febf9187fbed9bfbaf3fe3d2db4593b65602cf72a43765354df7a6bfba66b97b2f471fbadb656a847a7258f20e685bc81e55b243e9ad5c1ae8f41ef5ccfab4f6d14fe40e6e39a877b40b4a29baadd3f56de41c105fafffc349786cf0d2ec929ed2ccd3c296c1495c2db9c4f51873991782c91f80e68bd8dd30e8ea0aa0c45a9a9d0785c482001f9a978991c4cc92bd02c46243f3969447001b7aba89789fc55e9dc9936bcef0cb2e5d759dd2b29c0a2d537ec2de91c95e32d51d4944192669c8c896c782eafca17354222c230b24bbcfce00cb5190047e5c1dee1ed5b94c176a212888360a2fbb42feb0d26dcdfcd29524f7a565acc88ca10169fd34ea13ad4233cbf610bed13f1a3dbcaae6a707a9636a6d7e504501a2c8763100a30915ffb58ba9dcfad5d4f1253662e32a9c8ceff8226c7ae61b65cdb3a4309bdbf3431eaf58c34f2210df61291daa73325723965a0b1e379c97b6daab5d48835ff4682b30609fdc62a3aac9c0c07dbe3a1ef4e732e721f77e5cf72337c434a4786a2f974564e9321520bfa18cd42c21ef3dfba916bd99515ac37722449f6ae4cd14728fc48bd5b2fb45352df8d88a2a8eb0e3f39f2bf033d8d461b5a0510b245d6a8dd09c32c7fb08f72dacd80acbcfc2f1076ee22aae14c13da5d3f600eaec84c5e5506e3466309fafb98bb1a77f53751db5e2e6dc9dd4d042255e5e4133749e8d40261899c567aff6fc42276732e594fc336c01461f8e76770c7af52764416db3520b8f92cd7afcb2b0a72d25219a175bbad87b030b6e4746c264c6b51d55f72a686835ef92b255312463ac626bc06929bb985971a1941678127868282e67c4ccbd8c29ccc6fd8ee64f2ee7e69dfcac76f4c781e4ddfb6abc8ce9fcb888541aa81aa8d28c74cd95c125e38c0ba38ce96ba9a93be0027bdf6d21fca136fed96b5f7f8e0cc2b7346b303ab96c89fd839f0b88b95e31ccb234cf7631d31e288e012216b71f941536e331fb1386aea98d4ff0b930a17f265f2034c7380063697830be79a40ce4b3313e4f3917e26e4fea046430d6123553826f8bac301dc509ef2cf044ff4ef61f15034c980b7294aebea84d18c810a340d45fa6f9fa4dbcb13cfb9daceb01fc8fff87a09121f2316b13f30e8f51599c9f379646271e168e043280616318d6efc63771502b5424fa9e23f508b49edcf0e38cdad07847dd1a54244b563bc20da9fa43a71453e4b104baf0aaa5a033a484735e3315b129730cfed04089c12af0da83567ac3bae33242fd9a4104cbde141dd9cbddf104b14b9c822b817d06a261704af26ed55b09b58fa632294a6023ec6e1937beb962bd182d3bb1b446fd3513a29af0aaca9c30c049efa3c80e1c5aa41b3c942b29c6b462bc2cc0f3b31b3425120818c47f0b8972d8287b7d3fd601bcb9fc2ee9b6732777dde756007d27a5af56a1548364a11bc7740d068eba2156f58762112241e3f8fc8cbd564b4eed8ee20bec75204b8b78983d0cb092e38ca31720f8e821cb25f1c927189fc3919e945a466bf04b1fcc9300598e2e55f411bef2f0f631884cc0fcedad5e4eb0e98f99e07fa6c9c4c261354fbcaa4879c1d5ef20d65696508991edf642405780a64a090cdf407c86175d25ec5ce7aafbb1b258d3da745748c748783b315b256467b81a1ffb61bbe7b68b8252aea004a6ac07eacbc2947fbba31d90f97961586559b55cdf2d8605a26790e462dac063080bc10cc5cf84049b183e1852c27970ed5bc22f5a4b18ed8b408dc951d21a5858e579128e89381cee5aa217e7a956e24fcb2dc79f21e44a13bacd9bf7910ab4f6616ebdfd647aeca2c2459002eb744f15a53651690610468109b88bdcac44ffc70904b167957eda2c24e7f433633a3f7984ad9819960b166a7304a838e5578b870836f2e96b75566429b0bfd9b1f4f40fff4d8d3a28b9a0c662296b4d0543f345afc83c39e538be1ca0e0f0824727fc2ff13644cd5fe5f1eedf0ec0305904620b9f25e096d5ad045be85b8cb07cd72f337b2fc8e7478cf859a7b05d01fb9c96ab99fc877293570d3e669f6115ca4d297ad2488faef44840fc725693004fe4abfd76e9be3c2e58b06f1688b52261e58e0495c22d7dd5feb0f464353d5f9788488ddbb0dffeee33638d83ce8c420fb094f4c3c8212e84accc21965059ec30b4c920aa8b4c34b498e2397e88b88cab6a95431772d149b28bee22d6c1d924e9527f1b4c54712c508c2925902dfd5c1acfcb15277cdf31774fb74ade54c23bb9d839b228878348b3b7e06331c32d3f7aad137f004d0ffd0f48afb1b4ef5938afd353b2a1051b36d152f41e3950876ebc28881c30e98af4e1b7a7c4d4dbb1cc5682b30e1fdf55b4ab05cfed56eb0523967099e2f0041989decd7b3825e0ab6c0ab3098524ff3ca2af33e9efc6ef184530080acf04b58a1d30dd2f37f23df33cfbcfb5e0189b05bac5ed90df71470ddfa039dd5160579e362cdd5ef89b7041fc17017f9381c553184920ad80ea7c8aabfd0b9c0bffff43b4a38ebccd9bfec269245281b2f933d30d52d8c2f759f6fe2bd48b6098b4d83c7a44aed10aa1bfb0407154dad47ce3b1aeffd94dc14d73a19d3de6333e3879080c129b66b829d44c5d3e308ac13429be15047997f8009267be70f513142f7b260041a918af98a0d29d15c507c1bfd65f0e5bf6fd690785d2101de55c108bb2e4e699af6a35517c384981e694242111de41a128512279d6a630279b96c45602bbbd96d4d2895d3c45def19b07869b892e90187d2f0e01a0ef4db469dcd09e98fdc83b32c30797ef42b6e3b95c9da4a04231b015af22700a8c8840ba0ce4cae7dbffd24f73497705d5d0c4b273c7af173f1b7a1a6ac44d36fbc3061997ed5d37057cdac912dd044fab63d8bdce47af44305824688c18c7775ac5e7cc3ed7be5390660c171c931511ea107d904c21daa12f857c472ae8a25eb585e928368f79a2e3f21c355b5b18e6e7e6f1a5b9634b27d6501518c83170407900e9c66f013b33aefd09d96e3f174afc1a6cce995a0f0c52ec2295f34f6eca217d01f606207c794e5b4a8e17dfa1e950656febc2343855715bfca9938ab81da284b6deba93183d5af3f6e9eadc73ae645616ff55d72695030ae9d510f4eedbd640d2ece4e7dbf3183ef1483520b260467c29350f2c80fb15f7ce48a3c8284880e028bf4ac2ff395ff734d5f5105d3c5d02b3b614be189dabb566a36ac7e0ea0ec83693e303ac634737ec601e9a58665183a1e6e4ad5ab2448b9a02bef73d1c9fae2f38354d4a6d6a856bf6a812b5bd7f9cb05944714f558b1bb66d8d9fc398c53eb48ee238df9b989da08c8ad414ba3bc61db07192a62dfded1d97f1b42a87016ad3425322ba238096f0c0bde756d2cff26781b1f88814ff13dd4950a5cf69839aa81d8731ba04ce02f85eb6a5bba48c6be824afd01f98a1f64a08b0c19e54a26e4d8a966a001fd0cee38e0c673940b660f4e3da423c539da34fd167f13007ad8ff31d06d457394d92bb62a0716493601b85b820a6299a3d3798f411fcd7818fe9040a530f5169208ef2e774d7232c5cc4c563322f1b31ffc8ca18849876d0b8b4b2de84d7798d7a51a9a8641510f2e0fc571898de58f28dc4098ed877071c7f5d891c6bb29af1319af2e8edc07935aa4d876a66a2f2f14afdf62a66f7736617bcefbc7c61ec70f7ee8a41560779d559d3d42791c9071aa0013d9fbf88186a2dd18e02b9228e45305613a73f0e96373b5ba8993b8768d699ff1b8b786c15a2b2bed0747023119fca4387295b0a6fe5bc85652bca2ab47cbcbe248580ca690b4f230e278767bc45785a02718ac7501b22574c67049cea8dc2ac9c7b72a95b2846dcc8483f11975c06cc24db96c605f33afc3821f9cf5b0cb32f1f1df976e76cba121c12fb4850eaa1f4c69e822e863def50a935a345e592c5902931aebc970e96462d19f47aca01a3004f889936adee0ff0b62322af75a8c8b3a814e2713ede11ed443f932b4fae840778718eeb017bb5e3e617e887cf143fc25aed95e4a6b0d6119b5dba855a22b45878126a4f5691308d45aabd425cda09ac54f240d4d779ed8b8e2434d5f39a2e0956772eb737b813bd2bc8c52e4c0cf3ec52c575a207db69af71b9d343263ead0163f388fd2b5a999e397ac7829f985a10aa29abbc69affb07f6074f44e7ca209d451114dc5696e625d3b629fce09ad58520be0df5f57d8ac5d1a239b3f679f129fbad63fe364910a155d440a036a7ac1ab0bdf9cb03ed151bfc3b2c18aab5e4ae39945d3beb0631b418733888c4356e7c72', 'dce01cc72f1220b6dcd749ea6a939e1d'},
		ForsSignVerifyTest{'9f86d081884c7d659a2feaa0c55ad015a3bf4f1b2b0b822cd1', 'ffffffffffffffffffffffffffffffff', '00000000000000000000000000000000', '0543fb42fafbd65e1b76f99a8da5c7f0e9ee91975c55ef131865b1d024eed8181ebfd0a57ed329da90cfb63242df1b6c8eea72faaa484ea9a766e70219ff74bd4f7cfc769c08883102d365008b528291eb20d188e237328d266e1de65faf414eb7776847e5ddca12971cb8187952ea1196ee377971aaf7438baa5be231a93d78a83d0958750dc960bfe32f087b8b02d7124cd09083680007fe88f09f4ca6cb3e1fb14f81a6ffdc7c2d9852bf44787c0fea6582ae94fe08d40e5b9049716b3d3ff2e5d2776e4e78b7688e5a44be8bcfd7758b1188218db8471249e6271ff1f75b5fc0dd859db3491aee0f8dad52b1c9e48e31dfa56c9fb9b535110b42fd95f0d9dd8aa00c13737c61e6651a2330f46d47c4a0ccc873e87a4c918d0606971d95fd25be65f9be183e72cb0e720be5803ebcb966c7e6b0365f70d60bd19dfeffe3c8f0d960d523ad4ac8044dc1c451479623a617cfceae5da7a8dbd0e7e9aa3fe54505731faddbd094eeee36ec15ee168265e4894bd9ceeda29077fbba30e4048477aeac827bd6ff03f62b251dc05ca852f9c79f13276837d3315f923852aeb1b2d072a612d7d5198d1856ca5e621feaec924090a82cffaa671a497fd3074fc704b06d8bc0876e9080e1debd5a92b0d736c2af4a6d671bb7317c1d3313051aa72636c33a0c9e873dd51ceead201aade94a33339f96c2390e5bdf58ae88181c35040bf6f22e65c40a4da937a74eccd466e8451b144468e1790443c301412477062a71e7572cc290b5b3b0a36c0aa1cfd73bd55464e9b039965cfe0b3c1955d858e3ffa3027f1d113d88c7b46e42953e8be5b1a2e31b1b2db27029b849a3b6c1bd53e22d05a401914e8d8d695b02a076c1820f0b52781e7c33a9a2217fad4e1c930293293a71405d1bd4761489d2dee0613ed290ed5f4b5a1b69e657a190e8cd0af382845177bcc09b3c42136a4a7a94c5abf54a029497b1675b940bb2328bb645e7f39877d1526f7a95cf4b40924450c0bdc062cdaff598f63e164a6ecb28270d517422cae5be5bbb05e073947c632f290940a619a4b63be2461f7c4050117e903f00688648cbd3be4b5af747355d0c1e88725e5f35672931b8bad3fe63fe70a9b2a2c18893ef3089003114f5eb17a70fc533698766e6fff2b58cded815cbac258b249234e57130da085c5d488b9629ac829cc20f898aafc9deafa53833d840cce502d05f64bcf193e22a8539de576772591c113ef500f2ed31865321151e1c782223bb9139897aa87bfca221a983eba9db671aa4b1f1ccc6aadd9b57afc0e34fbb4a7253192b161e5d189fb608324808edb1181707dccbfff4e4228b5a028a3a9d8ffc2a3ca210fdda06007a710033433e859650a4e8df946b10c0af1fe77b0fc3695fdaff7b7128c4af666a70dd129bd647f50ea467e5a2c4ef858e9ef7c5f9fdbe32313f229515b20c31fe4d118090954bcfa60abdce2c4f03fecd4db5339293bec3de7b3bee82d41cfd79a8638201e61b5565cf3119b21d1f4fcc586c39e5617a2855ae1ab35c31259865ac9e070f70f12e36bff6eda66a16527aec28e1c1523e315aba44797d7fe300c0a5f1aab78dcbe449b7054c56ca75c37ed46e94cede204173210165cf9c16358423f84e8a8211da9c88ec0364e19ef7ffd0b472b72bb7476f30ef5b37f2cace531e238509c0b76ee7e47132d84856834cebeb440b7881f6b3c7f2c61a6e226deb9a32b5d3e7905e181ca91906cd4216acfbb28d481ca6fa3994ac8770aafacf693546839e545544ad187d214804012da8b94d1a72c199d414bd9bc49ca75ca0288405941d6f6ece34ae77b262c5a6428a5df705ff003382f14be993463a23de9e69a27c1324277fe675d92026c57cb099880413febe879733bc6918a6a62ab10b0c781d68ef6aa1cb61bd6be3efbd42fff1b417b4ffcb3ebcfc0eceaa3bd09134a326f6769840df0c7ae13719f36467522dc95fcafd4e1e0213c64a2615a2cfaafedde6b5b763d6019b15fed6a2460eda9ed021d710100251d53c7aefda71046c3c9971385755ef7dd6855f51e7ef5689eeba569b30c2510d7c26d52a8d7268b6d3b07002446385f356769c1fc1904e7a4ae6e7cb759f5fd280e7df74eae0a6cf67c7d650524a16b9e9b10e03546a3fe763e20b8fa2b5864c7d3fd9d1dbd1dc7867012c8d155987a27cbb5cb2d08af7d238aee50841b1afcb1821994461191a073c92bcabb3795e241e078b9eadc3c9ec5427f9b83a5e3ad5438c14db036c666ea18e44a36654826ee81b1c9215e61e08bc5d47289124e5d622b27a9a2e4fa6b35872315c5ae347daf346dfa4c2e43f770f36330b18b50df1cc5e081789312441ad2dab9dc3841f56a8d500db4031c6c8c1a301c246d610232222c5bd5e4fb45ac982735bf18db4881dbc6e0165cce6333655e181975b8fa601e9dc88c6a563638415d8fc4b28f8fd0c3292fb9b9600f443eebc6215b26d954bd70c7f481fa169b5ca6ee858b15388d070e67c38379616f40f5ddd9dd15ec7dec31e9f8b2a8b09cde6c4ca4dcaa8acc1a1f90b5dfb1a3580906b212da8304a9c3c019378bc2d4d0f35afae5a585a59091e1953150ef3819701dfa07dabdb7a66e5a644a5a5e9e5d7616b838c2726c830802b0fb02ba23e32fb2db603b53b5660d182bc4444bb52d435beeba4ca10d672cec880a27e1690b16be095cc74e84262023f84b1a7afaa2d0843d3eb4c2d45f377a4d3cb903058a8c11becb02b0de4af0e6284bc37f8d5bec0986ee355117f9037765425c9f05136f3781aae130639ada29f59aa2af6690e7fc0ac025a0d58205ded37e09b39339169430099556883bd1b8893996c41dbd110ff59e2f7e4f49c493383b20ba9b611aa9d5e6da282c3e03cdff65838debd61613fb616a3b80fd30ec5318cf55849a7575a60f2c5a374aa12d9bdf525bef466ca8edce0bec7a9e5d7081044ae89b1540d65e13436a3b8b985adbbb7d49fb3eb29ffb3c8389e57499bac2343d685a26d9061023eca34bc70f106c33e802b5785f8473fdeb612a930a9a96852a14145782876ffb0646625cdd97cfb535d4a6b5d3b1aeb0f99c4aae9e2d8634817f878b24b2a3cbdddbe4f782f024954f64d06b7b00ec8a6d6fa3788c63e7f8c1dcaec13f7844d78e37366a5ecc40f19bba5b1081892ea292674bb16f4f813c0d4f08f2ee40861ffb0cd6874a1ad8dd25f8d20119f6a362bdcd239a84c84233f254f944c62a9b0b79f0857fefd5984b085c92a2c7e66bf196c7718777e8fbace53a9621f33a3b0f7b4a2f2d48f136e8dde817036252f2bce5655ff51713b6d55b57be3263865783d0b69e899fd07f970f66c328cb51bc312753277bd4623f9f3eaecbddef0e3538477769e70098c42033daff1e33a41002d9310d476561bc7769aae20059f6463710fe2e0898ef685e0c338fdc6b350624aff7e95abeb4d4bb5d995f263983f05b242f7142ad5050f8ca0f1c1bbf26e066435f77384242b500ec7aff6d8c07ec43a16592307566b1ab295a1b815254684ee0e86dff080de5fa3e83ad1c1da7da5e188d7d4fbbe29619ef84d6058c5632584afab9a72105af416bd3727371de662de0c0d179bc57d2e71abbb7385fff3ad0e9af3d3897a8c7adf7992a7d786b33754d26ecb0287f9ea04a58c353c1286be080e07943e8233d964e137cad4f27e8979731381870d16cb0f3a9920a06424891a3e2a0775a1e673d70a4e63edb8a353c5677c3772d65350c3c3c71b95dfdb92bf112b0f62d578ecb4c91d3812ff35e7f24a9cfda52f04c09cb5d0a41e820fe006994868156fadf34e5b46f547fb89b8e3233db2d4facef4b369f951ce7e9a965e3c89b7240c20507a9e5cd6b07bc380325c820565bd03882dea434c63ce291f738a0958032c546ccaf05d3b6304df6a51d9f1300535f2e54e7a97de296191faf755af32ac5deec74c8eb02e9de0994fa3c77f232c96cdcd71fcfb5eb3357a7d8ccc69506cfb242e37888c057971dde92db6291789f2c7402747a6299417e07f7d75bdc1ba4184c6e68185af74dfed458a51cff0427dad4cff16a4c75db6714f92bfbc5fdc11c69977b098e4eabb5ab73fb3187252b337e2d667fa1308dd578ecf9c129896640fe1a1b3a3bbe8c480ce9f335b175918bd931928438348d53e32c0be7cfb671435f49247a645d4211c308674fcfcf9f7c9c0fad6bbcbde28c08e7b85561a6573fb604f9838bdea348d5ccaa76094e6e862419752ea5bff9f453c549674f872012f6d67b20973edc0b409904d3fea1362212554ca6eaa3fca3c4de6b9c5c11b0757f48dcecb3cbc134ae81dc9ee2fb0544df10ad1e44942eee5e4e50379fc4299b7d5355fbf4af432ff270f758b7e0d2fdcceb915c481ab7c678609e682acdab7c4d9a41590772bbeec0071ef83406459e96a9150fe6216c396c1a405ad3ac682b76edf7870cd9ea85d3f6f6b1cb70d18e51af707ef313acacb208409c6b2da04fc61b69bf89906564b48db8d8b7a537ebf3fa267d1d1cc8a14a0cf67559da939adff400f7af3690aaf9368edf34a723063a1dcaf01a5b3f32a6cb0828a78fa9c1034d2cacd95bc34bacb32f9247678808a8c81b5881f190bd6f14aec1ceddbf9ca562cc45788cd1cbbacfade21dc64b8416cab9730c1f5dd80e91279dc87df68f29253c10832e97e52479b2c7053a37f0ea728c820f2b2df8a65a9e79969348abd2fcd681cd3cfb4bf69dc86c747d8c2dbfefe281062e21631066d8ebaf68e448e92db116edd016f1fa58102cb2faca267ef1ddf64bbb6165cecb3772ce847983da8ced0be02c735886f4665e643b490b0d198d4e07e507d9b7b39a1e2f32e6b5f7b5e463e927055bef1c68c444246a84453af21778bf613a87e2f6d2d7d7f5c65b426444e02f6c7f315820d2f6dfc4163dac656a248e50a03aa526f9d9b3644196e526dbdd8c3b0aaf5c6549ce789a20caba74cb9f9b37152e2c879faa7b5586a9579398481b838288fd8aa982685569ca0f9713571698d24b3344e845d7fbe8a39f08c48930eff30c17d90cf5540bdc20bef2fe552ca657dbfe64673f2146ba9589baa5d8528d03d34a9bd44dc8bc282424392e27eab752ecf4b9556d3139ec17de3128a3ec30ec7039e6ad2106c31a3eb0846e3049c990611418477d9cdc9a479e315930f81022448ff5dc5964e1eb88951b24f0a8c1736149f49', '0bcbd03f9b6be9301cea5d617cf13a59'},
	]
	c := new_context(.shake_128f)
	mut adrs := new_address()
	adrs.set_type_and_clear(.fors_tree)
	adrs.set_tree_address(make_treeindex_from64(3))
	adrs.set_keypair_address(5)
	for item in tests {
		md := hex.decode(item.md)!
		skseed := hex.decode(item.skseed)!
		pkseed := hex.decode(item.pkseed)!
		expected_sign := hex.decode(item.expected_sign)!
		expected_pk := hex.decode(item.expected_pk)!

		// fors_sign(c &Context, md []u8, skseed []u8, pkseed []u8, mut addr Address) ![]u8 {
		sign := fors_sign(c, md, skseed, pkseed, mut adrs)!
		assert expected_sign == sign

		// fors_pkfromsig(c &Context, sigfors []u8, md []u8, pkseed []u8, mut addr Address) ![]u8 {
		pk := fors_pkfromsig(c, sign, md, pkseed, mut adrs)!

		assert expected_pk == pk
	}
}

// Test 3
fn test_for_known_answer_test() ! {
	c := new_context(.shake_128f)
	sk_seed := []u8{len: 16, init: 1}
	pk_seed := []u8{len: 16, init: 2}
	md := []u8{len: 25, init: 3}
	mut adrs := new_address()
	adrs.set_type_and_clear(.fors_tree)
	adrs.set_tree_address(make_treeindex_from64(3))
	adrs.set_keypair_address(5)
	sig := fors_sign(c, md, sk_seed, pk_seed, mut adrs)!
	expected := '2cac88fad4eeae791048fe07aa3544a9ab0db7949e4abe2d767811bce716bc008b512f3dc7992fe8d5fe70c0f822f65bc3c8f23ec667ac82a899d62267431e5957d9471da7421fc353f3a4e3117e5b826dbe311ae7149847237fcb470e4ca87ad9a1aac408b8b5e3083abdabbd7b43835cab0d526d48edb9394d2de1e336f032c927304c7d98006b391a246c026b4db4a7f9a4b9e23098d7979fa9e12596e91ed2e211744d165a6fa345a46f75466d7f9cf4246210a029514bacff2c5a7e388ed9367fb58b5e0822c3d626763ab284487c0ce3e00ef878da1eb86e79a644adb9a9594b1965a681ab3808b7449ccc3fad92c18b2dcf30f6039ba6bc905c0120c0007ee543f98332209796725f60c5215a9e22bbc28bc53a9ed7e80cd2b1a749ca15b17e02f21a655154fd0e376672843208e41bfcb86d13453a9acf9fa4fab1f9f0bbca7e8061a902626d4cf67daa1efdc250a680f1f7c73edd342e306fd5b6c583c863db88fc2ad9aa7cab71df150c808ee52368c247c00cdb6cd172148f621b05fb4c57760821ec6e0ff89b34a48d5070e9e31aace4ea4b3baab68d6fd8742629f156fd3f24cd7af90bd16bb7925ff6ae35d668a5fa16a6dccf53bb6a1fd84f43c6e5553c24889437ce33d1eaadcc7dd1a5725d47e1373d7b630afc3e6a4881f5884498333213de34b874f9e7156abe24df0d49ac1b47061682b1206adf3a90b7b187467375aa88e31b1998d2ca9ffb4f5b403cfa4986f058385d355d057049c1e39cba529da7ac0564d1042e7e19b91e45b9d93dcd7b47fe320e86065340aa02e982b098c7d4de76d35f90b49bc769f2fed7692d65bedd7e7faed34ac0d2b66e6cad8acb9c21403b6f188759e1624d7f3acc1475dc67b10120a9cdb61e5066ae48c47623acb8a22a1c448ae0a7526e8640c4c3c5fc39b102dcd5bf96e14a0cf92209e13e7de627d1dbc35efeec0adb0bededc8ce1e04726336114f8193fc22ed7c3fa25c57d2739e61c013a701e1f26b84e638d4a162a952da631b83ec82bd5c117842a1f3c90e4bd098c201ad01fa4826bb3f8f677f5a28bfb1341ae73830c2bde99049a98dd2e72203fe129ebb74df772dd23af9b65509ad64c9fe570c37a2dec3937d65a8742d15eb43232ade15770abf59f1d58dfb9e162288cb5704e575917584d91861d4d05c72802d8b0d20d60de536a559ec19863cf3df994f7f577e780d48fdc539505cf9cbe7d3366a98b19a3b4ff7c8ac873ba0fc7d8b62eb97dedc2b8fde1cd48769393c814858e26c5154a7a68f8fe04e89d51f2e9ea558ad893a93cf89c25e10560ecb52a1824a6950d9681113386ca46256d2f315196e491d7fddc302f2a6b13d209d01f1a931d73db8c7e526a3adb66374d421d2856bac4ae2273f5dbbfb41730e094037116e8c2c2142a2e99000a8651223be1d809f864dba1df1a351bd141e3823623b2ef41267c78b83d8348909e655ac0a6d7de7bc6869592c0c8098fdb0582d8d3f7b4b8d0cff1364c27ed916cc605ba0756c7de9547aeb18856b1a7ad47ab4216e65224064b781cdf331ec8b90069b8ca895711942ed015d94563e15cd15269691b2f5dadaa4de5fb65b446f56cdb15a56097a7ec21d2b8a383a5d57c9212d97ff49bda9e9fd7e4ac97a63a5d766b23951c46ae117ff035a8a01b6b13d552929030a39c93a6ce3514e849b9846d7cb50477d2f50c75defe9cf2e581aa6472c2d5091b174ea125546262026f88b809e883df0ca555542ccbf45463888eb69c4ae776d223fbc4aa9a3226a6902e08879e8f26cc5cc3c10e957b8b9df1d0f63ab2302d3848fa279887737582214fbaf2ca8c6d4db9a2dccbbf77436fc1c92094cc95f829c7d01537cf3e050db557f3af9f0666292566f866cf423ed7b3d319451f1c3a149fcdab3d0af11df4cea9f03091a50724d7e0828d959f75ee7a8dbd77173e0a8d9601d68359917b8322f1404d2df90bbbdff30cf95015991d269d8750342f87a9d128f71c1e2f59c4195c88568c33b2d9e3101c3d2eb8333dba37032ad1cecf93e1d9549eadcc51402b6facc0e9dc49eb319dd219e310d8685aad7eafa9eeb3c6a9ff8b0d92dd69ee21ae5ccba033aed106d353b3cf6f3ebc571bdd52d3564fae36fb72beb2c1e5560c10fc63bae4fd899e2477fc22f24f840bf707836ffc7555330a9d598529222e0a5236cd98a3fd7fe71397cfd5aadf18308e26952723ecf68fafef58ab686e103099877e3dcaf54017c3845037737dddc5cee97be961fc143c46c174debbe5dd50b54b78a6c3ed296e7ba807221df6f4edbcede1e112a8532ad4152a0451ee1ad5119f0b64febc9f70818fa91d3c20487846f6a4e0b6fdb58cd8c898b4674f89f58d340147da10af5534cc0a257f11ba2c56d5df3caf98dfe601bfbe5db517a4962ad1b5aef4e35fc09504564da0bcadff2a978c6bc5771db63afce16ca77afea52025207222936de1a4301b9c22cb7a82faae7e6de51c2a964ef6c5cd90f387438ada33d83d1298df59fc6655b89a44eeaa2193415d9a74288e1b938f7f8b3e3ff7b6cbd4dcaa4f94bdff08cc1d146be2b1b98288daee9465b9a559e0f45b3688a3e15d608625a605ab61c1ed68830af15af0a420a892b1a7d931398d38c693a682b831dcb2bd597cc6c688f6f8e1fef3af478e787b3fdcc973bfaec54bf35f95885f9dcbd4c2dec0e77685949e2e719f9efdcf87f68d53cc408a18cae49765c7e069db3589f8a40efd8079a2ce3d3f642ae810798ef005f164bc49a460f489fb6636de626cc9e15d9bac5b681a5778fcc47992067370685e2fe13fad1524b074ecc0c22b538f6a4dccc04e74bfeb8555e2ca70668e795891f2f29e90ee399860bbd304e4adc4b0fb906903cf76c14eae445f1264e9d02c9fdf8f136891a2edd673fd618fa9087cda3ee848ec664db24040ee9984b87b32f17426f874a1df9caf48e56189e7c77c5dcc7d67ae43ad8981090d194e7296ebe7fa4d2079e9459b3c94a9aea25417ea56c6b534a33f522e8a84dd72d36775098b0197bc35de831d4dd2e1b285ab3dc48f70e093b8e8371d163b4caa433b02300fa5c2e13151db1c007639f7fab7daddc7d61cecc434d98da5cd935bff6d6ff0249de2499f600247f45380421b8bca738f7706b3ac2eb72c0f063ec2fa49b4cd3eea81d78c05097af13e0627624f05b2a8ee35c1aee48d793d71376e520035a9adf3b4da3e5589fa9feb181e0760e42bebccc732d75278c8e3db0204ac4286dee76831debc5c747f739ce9ba8033c88395ec5c545f84e56b859af1e8ec8bed15ef95376dfd94080277f9a46c57be0d8dc95d8c081215984612108ce867d660219d82af26fc92ea0612984d54e2e9919ae21f9e707447b568fe377805ae91097130066735a71ffb3d2ee302a8238af655f78312a3114429d9229b70c0ca8a6b3610efdc3e255becaea51e210b3a953164461c2989ad008df28ee01894c6d004f3aff8330a0705e6dc310c114b507637df65ba9536eee7333a0aec3d066210876f18c68337e1c01557778babb9c42a3c22750062eb3d85f0b483d0df6fd1257ee50c51410c61bb736de6c5b299af5e1adea194a90b0df2141d4f09825ab4fb9b0677a81e0082b272d1d285de6f75d71be139e4c2600dea5382f25d6d31d2948fa2fb7b249f2c9d7d878b7d4fb83248ed9bf1d115f60790e04878b7aa6a06fc4777f6173167d6670f528654155181c837e1f3ce7a8878da886b2272edfecb480b011400d21e113516fb7e5ed586777c8b869b0daf770a8ee057a4ea9ec0c3e6173b569d4a9584d94154dd2dd398871e96fe74086565ad3de7f4082ac854cca03db02e1743a60610d0e9b280b4cf07324609d8a60696152e8a43e8d54dde2e4fa8520a2dfb1ad52e52b02d3a59f7efe0002fadb13cc4459a83adc9c95c7c629cffc49690e31e939838b10b099e6805e5f836afe87ddc555a60a170e420c4689602688e1bfdaf2acc8b8b7b5a2baa7fea26cee53a8234624f3bfa46b42de7e88b55be6b270673e514506dae3a3315721e12fcb6c9351840dc9190cc10a33b12a2c8458e2c7d604940278c225f4be63fb0aaa2b044cca2caa877f616ebc6c7c3d0925d8fcfa85ff9d7bb34cb583f67c2491404e360b8d44ba7bd5781212f14508b201ddec32f782a66f99524dc671dd9d6504b5157e05a9868de15601bac2adf0dd11a098641d2eb7e5e4bebcd0c0ac5bcd677ea268ab2e99bd60342400b5c212f627972cbe7131f09d96688254758bb15e0866aef3cf49d71e271bb5013e9678a2fe6b56dffc42f24fc8d3ffe2181c9396f84984be88f3fe6cb54876daa601e44294a340c52b64cd7e85b7a928639521f69ed9f62b2697d1a102f1f2dbd8ed8ac5f41c66206291fc7ded397c707edd225023323cc0065ea2d842feb8422e2c4cc91c7e0deb69e80cf3347a75585413fe33f6ec7be06ad09a68cc238b48cd58b8d4c900281b8cfa79d2afabeada78d80ff1c67844ad4277bf118864649a3ec6b28ae522ffd7533f98a5502b523d369a8a6a02de6f0840f44620f206a48b6ebd0120e8e7f311e3b61f09a57f499c6931d475021bb9637ce37c0e657720e2fc2c04595a360725575c7f9e90eb41dee5254476d1fba11f3c19b4ade31e888e919d3f30030f3a19605154fa89d14f5fe7d1c787aac421f5c3ddd3b69f0a335c5605ab674f705305b0a5bbebf4202cc5023b47b21eef6815e0f6b08d2b2da46323938729bdd55f5341ff14d36df69803229c6046b2503a62d4e47da0195d0028cbfe0a67bf5230b4b8a8d2c1c31203ceac2873a860c2355e5f859a2be634f323dc30efe4ce3ffa7a61e0a32ca8d3a4cc611bee7c0f08ae0e7c17c2a9c8e42d5dc22e315b39800c435391233c937ed90125ffc463573afb4c15b452d653e03de6b13497a3e6e2757e7f218b4b8c0430d9a27c26997b092f20985c4af70d1cf2fd0d42d86732d80711fb25ce2e0a2a1ae179073350832cf4495ec887a77739598aabd4f3caf2a2c70b70631e0fe67e3ee4aa7843c41c2f253bc696d6b859844e28f9a416314a1d740cb5e757000ff1ca5422dafc98a3cd856ee679d11f9d4fe0ff7f1e6e9217f53e74bacc9f8098d1c7e54e9ed32f69f06e2b5a345df79c4d3864078ec89befb5585cdc3d79e51bd5fe70896089ea2af20e99b6ca2ce814190f602542a1bfa738ea'
	assert expected == sig.hex()
}
