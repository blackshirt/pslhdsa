module pslhdsa

import encoding.hex

struct KeygenTest {
	tcid    int
	kind    string
	sk_seed string
	sk_prf  string
	pk_seed string

	sk_out string
	pk_out string
}

fn test_basic_slh_keygen_internal() ! {
	// slh_keygen_internal(c Context, sk_seed []u8, sk_prf []u8, pk_seed []u8) !(Sk, Pk)
	for item in keygen_samples {
		kind := kind_from_longname(item.kind)!
		c := new_context(kind)
		// dump(c.is_shake())
		sk_seed := hex.decode(item.sk_seed)!
		sk_prf := hex.decode(item.sk_prf)!
		pk_seed := hex.decode(item.pk_seed)!

		sk_out := hex.decode(item.sk_out)!
		pk_out := hex.decode(item.pk_out)!

		// splitted from pk_out, where its pk_seed+pk_root
		pk_root := pk_out[c.n..]

		sk, pk := slh_keygen_internal(c, sk_seed, sk_prf, pk_seed)!

		assert sk.pk.root == pk_root
		assert pk.bytes() == pk_out
	}
}

const keygen_samples = [
	KeygenTest{
		tcid:    1
		kind:    'SLH-DSA-SHA2-128s'
		sk_seed: 'AC379F047FAAB2004F3AE32350AC9A3D'
		sk_prf:  '829FFF0AA59E956A87F3971C4D58E710'
		pk_seed: '0566D240CC519834322EAFBCC73C79F5'
		sk_out:  'AC379F047FAAB2004F3AE32350AC9A3D829FFF0AA59E956A87F3971C4D58E7100566D240CC519834322EAFBCC73C79F5A4B84F02E8BF0CBD54017B2D3C494B57'
		pk_out:  '0566D240CC519834322EAFBCC73C79F5A4B84F02E8BF0CBD54017B2D3C494B57'
	},
	KeygenTest{
		tcid:    2
		kind:    'SLH-DSA-SHA2-128s'
		sk_seed: '20D43B51FB11AF1FE3C6459B7BB90D50'
		sk_prf:  '4F63BA1D6CC9B355D47E49C958658160'
		pk_seed: 'F420447CFE8F1823CE5BBFF0030CC69D'
		sk_out:  '20D43B51FB11AF1FE3C6459B7BB90D504F63BA1D6CC9B355D47E49C958658160F420447CFE8F1823CE5BBFF0030CC69D31A2F32390C22B1AB974B5F5A2B3844E'
		pk_out:  'F420447CFE8F1823CE5BBFF0030CC69D31A2F32390C22B1AB974B5F5A2B3844E'
	},
	KeygenTest{
		tcid:    3
		kind:    'SLH-DSA-SHA2-128s'
		sk_seed: '94FDCD4EDA1BBF7FB510FE16C42BFC57'
		sk_prf:  '2859455BDA66A81FE212501B3D82572B'
		pk_seed: '357DBB62C05296027861917D4AA53CF7'
		sk_out:  '94FDCD4EDA1BBF7FB510FE16C42BFC572859455BDA66A81FE212501B3D82572B357DBB62C05296027861917D4AA53CF7DF891E96BA5C7997319F7D39B2B455D4'
		pk_out:  '357DBB62C05296027861917D4AA53CF7DF891E96BA5C7997319F7D39B2B455D4'
	},
	KeygenTest{
		tcid:    11
		kind:    'SLH-DSA-SHAKE-128s'
		sk_seed: '2A2CCF3CD8F9F86E131BE654CFF6C0B4'
		sk_prf:  'FDFCEB1AA2F0BA2C3C1388194F6116C7'
		pk_seed: '890CC7F4A46FE6C34D3F26A62FF962E1'
		sk_out:  '2A2CCF3CD8F9F86E131BE654CFF6C0B4FDFCEB1AA2F0BA2C3C1388194F6116C7890CC7F4A46FE6C34D3F26A62FF962E1E8C88D2BDCBA6F66E50403E77FA92EFE'
		pk_out:  '890CC7F4A46FE6C34D3F26A62FF962E1E8C88D2BDCBA6F66E50403E77FA92EFE'
	},
	KeygenTest{
		tcid:    12
		kind:    'SLH-DSA-SHAKE-128s'
		sk_seed: '35DE5545D627E5AFC8F8669662A8728C'
		sk_prf:  '51569550F70E010898462443C877CAAA'
		pk_seed: 'E756D06936FD4C3B6E41C5013D2B36BC'
		sk_out:  '35DE5545D627E5AFC8F8669662A8728C51569550F70E010898462443C877CAAAE756D06936FD4C3B6E41C5013D2B36BC44C0B9567B59F7A02D3034CAA491129C'
		pk_out:  'E756D06936FD4C3B6E41C5013D2B36BC44C0B9567B59F7A02D3034CAA491129C'
	},
	KeygenTest{
		tcid:    13
		kind:    'SLH-DSA-SHAKE-128s'
		sk_seed: '47098E209EADC5C15FEC2B2E58F3016A'
		sk_prf:  '9B9054CADFB443724F253FAA7F2178BE'
		pk_seed: 'D4CAD475F7579DD5E29562F962188C27'
		sk_out:  '47098E209EADC5C15FEC2B2E58F3016A9B9054CADFB443724F253FAA7F2178BED4CAD475F7579DD5E29562F962188C275D0AF4241F0F622E05BD10DA0B70B3FB'
		pk_out:  'D4CAD475F7579DD5E29562F962188C275D0AF4241F0F622E05BD10DA0B70B3FB'
	},
	KeygenTest{
		tcid:    21
		kind:    'SLH-DSA-SHA2-128f'
		sk_seed: 'AED6F6F5C5408BBFFA1136BC9049A701'
		sk_prf:  '4D4CE0711E176A0C8A023508A692C207'
		pk_seed: '74D98D5000AF53B98F36389A1292BED3'
		sk_out:  'AED6F6F5C5408BBFFA1136BC9049A7014D4CE0711E176A0C8A023508A692C20774D98D5000AF53B98F36389A1292BED3F4A650C56C426FCFDB88E3355459440C'
		pk_out:  '74D98D5000AF53B98F36389A1292BED3F4A650C56C426FCFDB88E3355459440C'
	},
	KeygenTest{
		tcid:    22
		kind:    'SLH-DSA-SHA2-128f'
		sk_seed: '70B19FCA9B6522347E32344FF3293053'
		sk_prf:  'B4ED68C937BBEAE268A4948C72B044BA'
		pk_seed: 'C5BF30C4A6787951315A0126C16566C9'
		sk_out:  '70B19FCA9B6522347E32344FF3293053B4ED68C937BBEAE268A4948C72B044BAC5BF30C4A6787951315A0126C16566C9B2A4A872833E75A686AE7371F74286B8'
		pk_out:  'C5BF30C4A6787951315A0126C16566C9B2A4A872833E75A686AE7371F74286B8'
	},
	KeygenTest{
		tcid:    23
		kind:    'SLH-DSA-SHA2-128f'
		sk_seed: '35C317B8625A0AE432CAA14D3CACCB90'
		sk_prf:  'B0144CF517FB109EBC880DC8361D1CA6'
		pk_seed: 'D7036D522C1FE1CD6EEA07DE0ED5D657'
		sk_out:  '35C317B8625A0AE432CAA14D3CACCB90B0144CF517FB109EBC880DC8361D1CA6D7036D522C1FE1CD6EEA07DE0ED5D657C497573D5093F4AC806142A550F30621'
		pk_out:  'D7036D522C1FE1CD6EEA07DE0ED5D657C497573D5093F4AC806142A550F30621'
	},
	KeygenTest{
		tcid:    41
		kind:    'SLH-DSA-SHA2-192s'
		sk_seed: '3BFAED208B7DC795BF3647F86E4B48BF9ADB8D6784C50155'
		sk_prf:  'A20311739497C3FCB860EE47E09EDE036F7AE8A939155BC0'
		pk_seed: 'A67856A81A6ADBCED7F1A2780CC48A06681BA5E8C7938506'
		sk_out:  '3BFAED208B7DC795BF3647F86E4B48BF9ADB8D6784C50155A20311739497C3FCB860EE47E09EDE036F7AE8A939155BC0A67856A81A6ADBCED7F1A2780CC48A06681BA5E8C7938506BD031BC8124F95F0BAE2BECB2A3FBBAEC453C04A6E918FFB'
		pk_out:  'A67856A81A6ADBCED7F1A2780CC48A06681BA5E8C7938506BD031BC8124F95F0BAE2BECB2A3FBBAEC453C04A6E918FFB'
	},
	KeygenTest{
		tcid:    42
		kind:    'SLH-DSA-SHA2-192s'
		sk_seed: 'A083FDD6DAF6FBFC82F879F69AA2B9AD2B7C722585B67598'
		sk_prf:  '4A57A583ED81CDE66ED87634A40A67AD64486E19338C13D7'
		pk_seed: '854D536E8EEC3E703E1248E611AE16F29AB332D1F8A7EDED'
		sk_out:  'A083FDD6DAF6FBFC82F879F69AA2B9AD2B7C722585B675984A57A583ED81CDE66ED87634A40A67AD64486E19338C13D7854D536E8EEC3E703E1248E611AE16F29AB332D1F8A7EDED57D6FB440CD07BEAB081A4F6E3D003262DB8CE1931EB60CD'
		pk_out:  '854D536E8EEC3E703E1248E611AE16F29AB332D1F8A7EDED57D6FB440CD07BEAB081A4F6E3D003262DB8CE1931EB60CD'
	},
	KeygenTest{
		tcid:    43
		kind:    'SLH-DSA-SHA2-192s'
		sk_seed: '72D9AC9CDCD347FA90479F908A4AFA7CA972DBCF0BF2A5DF'
		sk_prf:  '760555465A27F5B47B43EF53C6EC6441B8C2DBAD7FAB3C94'
		pk_seed: '0A3D81B32C499138A1FCF22F927680CB33E3ADFED3FAA546'
		sk_out:  '72D9AC9CDCD347FA90479F908A4AFA7CA972DBCF0BF2A5DF760555465A27F5B47B43EF53C6EC6441B8C2DBAD7FAB3C940A3D81B32C499138A1FCF22F927680CB33E3ADFED3FAA5468AE272BB8AF09A3445A3F3E8F9FB70B6E20BDE23C08C75F6'
		pk_out:  '0A3D81B32C499138A1FCF22F927680CB33E3ADFED3FAA5468AE272BB8AF09A3445A3F3E8F9FB70B6E20BDE23C08C75F6'
	},
	KeygenTest{
		tcid:    61
		kind:    'SLH-DSA-SHA2-192f'
		sk_seed: '45D7131C727DF1CC51DB85B44E37868215DF8AEC5D1B552F'
		sk_prf:  '92BC5FC8A2969FE0A522492082E994DE1DDC90FA984F847B'
		pk_seed: '8330589C20701AA9F11B473B67E1D67E1C6A2EB6C86265ED'
		sk_out:  '45D7131C727DF1CC51DB85B44E37868215DF8AEC5D1B552F92BC5FC8A2969FE0A522492082E994DE1DDC90FA984F847B8330589C20701AA9F11B473B67E1D67E1C6A2EB6C86265ED13A3EA895C4EEEADDE8A796BBA5233F0D86EE5CBF2A6F99C'
		pk_out:  '8330589C20701AA9F11B473B67E1D67E1C6A2EB6C86265ED13A3EA895C4EEEADDE8A796BBA5233F0D86EE5CBF2A6F99C'
	},
	KeygenTest{
		tcid:    62
		kind:    'SLH-DSA-SHA2-192f'
		sk_seed: 'C359F4AA77D938A79B7269C591A5D8120F882F00932CB633'
		sk_prf:  '6715B05D2B057DD0E3822C5E316D25381D85591F37EA21E7'
		pk_seed: '7B3C40FBA0598852B9EF5045DFAC695D3E69AA20106F13F4'
		sk_out:  'C359F4AA77D938A79B7269C591A5D8120F882F00932CB6336715B05D2B057DD0E3822C5E316D25381D85591F37EA21E77B3C40FBA0598852B9EF5045DFAC695D3E69AA20106F13F4CB7B1DDBFB5D8623004CBCE479DB132A48DD47C4F5171E16'
		pk_out:  '7B3C40FBA0598852B9EF5045DFAC695D3E69AA20106F13F4CB7B1DDBFB5D8623004CBCE479DB132A48DD47C4F5171E16'
	},
	KeygenTest{
		tcid:    63
		kind:    'SLH-DSA-SHA2-192f'
		sk_seed: '809EA380F5D42FBC8DFC75E90C42820B37652EEF2CA7F5B6'
		sk_prf:  'DDCFE30EC2D375032F4F3C032A5AF4D6B46C7556D5D84B8D'
		pk_seed: '808AD21AF4358E1696E09055A39F265712FA466CCCE4CB8B'
		sk_out:  '809EA380F5D42FBC8DFC75E90C42820B37652EEF2CA7F5B6DDCFE30EC2D375032F4F3C032A5AF4D6B46C7556D5D84B8D808AD21AF4358E1696E09055A39F265712FA466CCCE4CB8BC33F99596B2009A4956E0318F81FBC63A69D0FD1BD96F04D'
		pk_out:  '808AD21AF4358E1696E09055A39F265712FA466CCCE4CB8BC33F99596B2009A4956E0318F81FBC63A69D0FD1BD96F04D'
	},
	KeygenTest{
		tcid:    64
		kind:    'SLH-DSA-SHA2-192f'
		sk_seed: '411191D5555C3C1BADA4F81EE616E79158211EAF57D29702'
		sk_prf:  'E14A4DE287CD88FA06F29B8E6BF33AC6AFF7245938585B62'
		pk_seed: '801E3905E31F66F06DFEE8C553F49185717DB104BA382893'
		sk_out:  '411191D5555C3C1BADA4F81EE616E79158211EAF57D29702E14A4DE287CD88FA06F29B8E6BF33AC6AFF7245938585B62801E3905E31F66F06DFEE8C553F49185717DB104BA382893AE7B7E408E80A4A0488FCCB6D137DFAAAB7328DED1DFF3F0'
		pk_out:  '801E3905E31F66F06DFEE8C553F49185717DB104BA382893AE7B7E408E80A4A0488FCCB6D137DFAAAB7328DED1DFF3F0'
	},
	KeygenTest{
		tcid:    81
		kind:    'SLH-DSA-SHA2-256s'
		sk_seed: '2FBEAB9A6A80FD817E7EFCDF834EFBD4F0A36195D7598408A6A151E93DE6A557'
		sk_prf:  '5D0B37D1ECBC68265B0AFEECBBA783DD27EAFDBDF3143E4AF3E5057FD5C2DADA'
		pk_seed: '1322F94917AE67D0DB420203178D591283C08BE8A1385A16CE70CD9FBAFD2AC6'
		sk_out:  '2FBEAB9A6A80FD817E7EFCDF834EFBD4F0A36195D7598408A6A151E93DE6A5575D0B37D1ECBC68265B0AFEECBBA783DD27EAFDBDF3143E4AF3E5057FD5C2DADA1322F94917AE67D0DB420203178D591283C08BE8A1385A16CE70CD9FBAFD2AC640041EAB68A4A653F89CAB7585F6B410603326DBBAAF733E7E72CB6097A4A452'
		pk_out:  '1322F94917AE67D0DB420203178D591283C08BE8A1385A16CE70CD9FBAFD2AC640041EAB68A4A653F89CAB7585F6B410603326DBBAAF733E7E72CB6097A4A452'
	},
	KeygenTest{
		tcid:    82
		kind:    'SLH-DSA-SHA2-256s'
		sk_seed: '59DC672E7B975F8911409FA7FDE582BD14AB3CEC31A57710155E8AC44C5A5649'
		sk_prf:  'A9E7E3F364C34815AAD9215382250ABBB381CD424E43DF32FBAC3056AE71B809'
		pk_seed: '4F08486D0D98C7DEE706594123BFE3DEBBCFF15BC7CAEAD58DBEFCCB34274B9A'
		sk_out:  '59DC672E7B975F8911409FA7FDE582BD14AB3CEC31A57710155E8AC44C5A5649A9E7E3F364C34815AAD9215382250ABBB381CD424E43DF32FBAC3056AE71B8094F08486D0D98C7DEE706594123BFE3DEBBCFF15BC7CAEAD58DBEFCCB34274B9A6483E64DBF92D7332E2F0492EBD21F3935500E450F45DEF5EA588C2433F6663B'
		pk_out:  '4F08486D0D98C7DEE706594123BFE3DEBBCFF15BC7CAEAD58DBEFCCB34274B9A6483E64DBF92D7332E2F0492EBD21F3935500E450F45DEF5EA588C2433F6663B'
	},
	KeygenTest{
		tcid:    83
		kind:    'SLH-DSA-SHA2-256s'
		sk_seed: 'C5C3D80CB42286F9C24BB078D3FAB98093B9EFE0083835373F2C7F85A7275704'
		sk_prf:  '5E33775CFEAE650C53926A86F9ACB5D749C0F3B9FA5B37534CAE3C86A7CFEF67'
		pk_seed: 'DBEFAF8E209A7B5DFD3FC92C56DDD9C505085054417FAE0A440D121FF1A07371'
		sk_out:  'C5C3D80CB42286F9C24BB078D3FAB98093B9EFE0083835373F2C7F85A72757045E33775CFEAE650C53926A86F9ACB5D749C0F3B9FA5B37534CAE3C86A7CFEF67DBEFAF8E209A7B5DFD3FC92C56DDD9C505085054417FAE0A440D121FF1A0737130ECD796BBAA118148425CB8493A57052574862806D56A0BAEE6F1789525FB06'
		pk_out:  'DBEFAF8E209A7B5DFD3FC92C56DDD9C505085054417FAE0A440D121FF1A0737130ECD796BBAA118148425CB8493A57052574862806D56A0BAEE6F1789525FB06'
	},
	KeygenTest{
		tcid:    101
		kind:    'SLH-DSA-SHA2-256f'
		sk_seed: 'B8ABC485122BE003CF36D677BEE7F47EA1017C39D96D0C56A87A7ADAD24F731A'
		sk_prf:  '9222684FFACF803D44CB98222C44B3C519698B798D8F7A759FE2FA6EF173CF64'
		pk_seed: '0D50E82BEDB42E03CC967E7FD24C12777855A946FD49471184330F096A75B561'
		sk_out:  'B8ABC485122BE003CF36D677BEE7F47EA1017C39D96D0C56A87A7ADAD24F731A9222684FFACF803D44CB98222C44B3C519698B798D8F7A759FE2FA6EF173CF640D50E82BEDB42E03CC967E7FD24C12777855A946FD49471184330F096A75B5617FB65FBD08D05F24F20CB3875E28FAC4A52A2513C7EF447B8E9328632A684CF7'
		pk_out:  '0D50E82BEDB42E03CC967E7FD24C12777855A946FD49471184330F096A75B5617FB65FBD08D05F24F20CB3875E28FAC4A52A2513C7EF447B8E9328632A684CF7'
	},
	KeygenTest{
		tcid:    102
		kind:    'SLH-DSA-SHA2-256f'
		sk_seed: 'EFBF2801445EA159BFF2C460A3A09FB03C5E47547C9621A97B1CFDB7B265EBBE'
		sk_prf:  '8079D79F1559A5F9FA2D75C7C2D0CEA6A531968EE97AB4B28EEFE8A11D685E86'
		pk_seed: 'DAEFD98FFB246D311128FD58339EB970C2310849ACF011AFC79A40DEF5F6A661'
		sk_out:  'EFBF2801445EA159BFF2C460A3A09FB03C5E47547C9621A97B1CFDB7B265EBBE8079D79F1559A5F9FA2D75C7C2D0CEA6A531968EE97AB4B28EEFE8A11D685E86DAEFD98FFB246D311128FD58339EB970C2310849ACF011AFC79A40DEF5F6A6615403936464A0CF48C8FF5AE356A1ADEF9B4245FBCE06BD4918A442300E3B12E7'
		pk_out:  'DAEFD98FFB246D311128FD58339EB970C2310849ACF011AFC79A40DEF5F6A6615403936464A0CF48C8FF5AE356A1ADEF9B4245FBCE06BD4918A442300E3B12E7'
	},
	KeygenTest{
		tcid:    103
		kind:    'SLH-DSA-SHA2-256f'
		sk_seed: '35925CD7C6F00268C3F9481D03D8B9504C249647BD93A4ACCB0D44D404F54657'
		sk_prf:  '4FF44753D29B314C0EFFF3C14E3B23E69BB96F25596411604B25215AC4C8FFEA'
		pk_seed: '19F753852878B9FFF6734321B3DF5548F89D9FE40CA38D942EF25FCD48D35E12'
		sk_out:  '35925CD7C6F00268C3F9481D03D8B9504C249647BD93A4ACCB0D44D404F546574FF44753D29B314C0EFFF3C14E3B23E69BB96F25596411604B25215AC4C8FFEA19F753852878B9FFF6734321B3DF5548F89D9FE40CA38D942EF25FCD48D35E12B090FD27D955951A4199F0213A0F95E488ABC48C2B99F1C5112B4AEBF3A246B0'
		pk_out:  '19F753852878B9FFF6734321B3DF5548F89D9FE40CA38D942EF25FCD48D35E12B090FD27D955951A4199F0213A0F95E488ABC48C2B99F1C5112B4AEBF3A246B0'
	},
]
