// Copyright © 2024 blackshirt.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
//
// The main SLH-DSA Signature signing testing module
module pslhdsa

import encoding.hex

// Test 1
// Test basic signing and verification
fn test_sign_verify_internal_basic() ! {
	sk := slh_keygen(new_context(.sha2_128f))!
	pk := sk.pubkey()

	msg := 'hello'.bytes()
	addrnd := []u8{len: 12, init: 0x0f}
	sig := slh_sign_internal(msg, sk, addrnd)!

	verified := slh_verify_internal(msg, sig, pk)!
	assert verified // NEED TO BE TRUE
}

// Test 2
struct SignShake128fTest {
	sk        string
	pk        string
	message   string
	context   string
	signature string
}

// The test material was adapted from golang version of slh-dsa
fn test_deterministic_sign_verify_shake128f() ! {
	item := SignShake128fTest{
		sk:        '6c1f4a3889984abd0d30e9454e8ae15d423be3aa1b0024599639b0bfb9c41e9fff34692100a04a8e9bea7ab80e2eaf8031e099f8dbdd09e71adf94836e3350b1'
		pk:        'ff34692100a04a8e9bea7ab80e2eaf8031e099f8dbdd09e71adf94836e3350b1'
		message:   '74657374206d657373616765'
		context:   '7465737420636f6e74657874'
		signature: 'fe9a71dc6a6920b113a168b78fdf75e0c33edb3d7302227abc8ed4c4c71def4b2b1ed071eb57129ab6387b43e2ddd659454eb1039fbc61b00dcdc0babaa844bad98628ccc862de4e969b6457ff21fd4cf538a50b89e4b7d77a1554ba16137a4c566e0e5d450876f2dfc4f90b18a578cffeaaad93064f8a5bed56e6a5d98e477253c133899c42eec2896e025f3fffe92f5148ef7875345c223f4fe8a6bad0a50717553037e103acf0d12d0dfd3fa71d30ca2bbc0253ce4d01fbad2002dac53fa029e2c0cc9e9f551e737646d63921aed8558862005b06793a8ebbcb099cfdd83827a4314ec6587485ecc3d93062e93be2d78039e6ca9bc03b12c1562fee0bd2e5cdc7a5614922b8f9bad9ae65f8889db82ae7f5ecb67c34289eed5c34abc8784b797725c07b219dc54cd9991031cd802b84c2b9e0429feff755c1ab380d79e0c7f7bec55db87d5c18517d75f0b2866da80f6b61b07f7394c56486ba1e1da16798f909441158e2589afb2f72a23321e793266573e1328d11fc26ca792de5402e1f6de8615832344a7779f72555448e3ad3795cf448d09d74ba56de6c364f14a6ea3cbacbbdc2a41751e0d213859f9f74e3a78e98afc4df9a04eee68fe86031c101ed43dc32d9ddb85011c04cddd298134faef2c11e0aece865f497c88335741e8a85e5866c2473eb27f9c9a090e79ab49dada78fca2faf3a85b2572a5866ae4ff224c8451920198c04a5d984caf225efce8bbab7dd7967a2719bf22f89529deeb38fb8f880cfb2fd2d2ce3f7ae433260f7bdb78ad78d4f3f506d07a4febf95a7b5ad431081c88b030e9869107a6eb5526c871eae188bbb6428e067150d504ed508b3bf11f0e61f01b11ec0ab26de6e75cfc2ab92b7fea9d3763b4bea54c984c18daa5a3974d9bb93454a318a9193e9e1cf7d24679449dc2d40b11fbdb58bd46c4e3e572b6bde4380570c58fbb12d4bb7c2fb60a7911e8d336e16c55d56c083f69c64de8ec1bcc4bb1b2d09d8af9de23ff6c39ca53471e93f152bc5e51d59edbd6e5546666519f5153e3efe621717c42c96a20876eccd3f93f7a82fbf6595a7af2a57754762bbd31936db4c77d54362d15f37eb7cd72e7ddd940792b3992bff15f81c28a8b1dafa34e217b5bb407f9f16fe2363cd8f063f8548b35cb123d06615133f1672448bc3131b7c5dd5607975dd3960925fa02e984ab4df6cca56b5e24f1b5939621b7777fc919168948769eb912fa160ec1cfbe8284b4c57a59bd9921bb0666a95d5379f59a70b8d232e5c055d9251a90029b9a8cb75a32f54297ae5b4d0c0e7bfdd2a202d65dd52052efa43f60c795c898ac8e6852caba5a8304cc814af44a8bfc97e59043d2487a9724a7a209feddb490ddf17cdc5ea58fa4759e912adcddfc0c43b8a050fd143a2dfdc7f4f9293630792455a03af832212cf82bec2979c89887da4f5f211e8638b7b6eeaf5ea4a22cc72fcd83629215a325f4930027e6584db476269ad47da2948ea3ca87e856a442cb2a4bef2b59b208965d4c5bedb3d8bd10a608b13ef1eb9c06438a2a16b8fe6ea9e35cc346591e3199de6581b5cf81883f82a010614cf52579823a802d2981ee13689b3b29412133a6b7c18030007da842af81f510754468fe90b0b2a2dff44a186104669432dd793bae29ea1793966c43438d4b190d414ccd0d4455c837c55d694308dfd53403bb0cc4b255f56d9329cab21ad44a72f5e5d02fa939c59b5787f3ccd503e95eaa8141387b6d55ea6fd87b519f8caa146a4e60a7071645f3344a3b1af79c4f28367c9120738b4d91945899d958353be4a84a73849e268399a905202e5e3947fde7aa7fd7266222f579a1140f4b5f412b18a7c6e6404eaca3eca437d2bd9723f405eb4f36947539696e6e0901475c99e26b540a3845101125dc1f6d9673d432a48b70344dda574b155c6fc098d241b657c508b45e6a0ea7d8cc79e80fa03f0d24452c63b4bfa90db6e85dbd38c5fd7c09236a8f20a46045216907a14743e638afe760de17542d6d4b2bd121ac1aeb836d3642f403998beb65f865ab9a6fcaa6d0906be63ff0e6b15f387e5c5ceff8ea4d23e06491bdf7dfe3d24264ae9afdc3e25ac8b3362a2c2c4e0ae9fbdabb209f4b04371912864d486a6a000a88ebea1e01b8a6ce96af157fbb8393672d0b8d9e629f9c6c40145ec66dd118a56805919aff3aa96dacd44a3a2bf9160b28ad15fc69ef89da0116a514f05a72a9b98811f6fc9b08214464e3d053a92fad9b7c3a2b9ba10301a81b561c7028f61e222cd2da7e87abd4196b0ac45706d62400fb2c8f0f9b153ccdbc47ac6f0c74d50e276c3820b40355ce90800692b700c59dfce9a410279bf63c29ddf9e673a36e199804e64ac1f494b8e65a1403da48acae189fd4685a245da10d41786234f3b12a11d7e3dd432ba1ad3f084cf45eeeec8a3b5d8991110a34949eb861118d25e3f06c0032bb233da15004db519042e62c359401c7e832534dd912d8b261ae255a5390d85f40bc4e3ecd4eef091aeb9b15b5f4f0c0e02d2c00db095e3c5d3c57275e45ea41d37fcab6f04d807ca96c90c26d7d0c7c2d691dc1870944d9226ff8efa143bc8d48be6ff438e951d21841df58f91fde297b07cba4b193c6d93aa92a4044e886bcaf4bdaf7b3dddb80f348018c9e55fcda8d86372b0da9d219034b635aaf15d711b62ce4bbe30a8216239f80db0a9ab3bdfd6e2f022c36798d72ef6467731a657d5e511c3234f9dfa6db158506f5599eb82dcb79375caea8ce3e786a901bf791602ecef231dcc07a7ed34d346e8581b5dbea796e70bad5c25135a73d1e89b4264f7333a2859b348261d19cdd0b1c6d7aa5cb65d79dbd6618f1fa11a65621af049a30c855066385c4632f9f51b3b4aed9107f395da9adc3bcd2b0c19a6d0ddb1835616a5cc97a1d31d25b8dcdfb68956d79120129c31c3486258ab7d8e36f15581d1138831a5d6be2dbaeeb9c9dcf7b86fa16a75902658650a6c5e81b400dad0666efbd04c2de45b910e73eef4669a142999cc6aa4bb79666b8ec686a38a85be7bcecf9de5580c78b621f752eb7b0e1dd11348d4f4024f3383121c968fc8fc05d692c2dc586b3c0dc47246143cbcdee6a1fa16552decb60466b40dfedb44133673fabc16d8466a7289db3cd5132b3bd14979d5ae8dc8ac54c6d759d608236721cf0deb8b9f73d68f77f58e39b41c351f32eef7d5804695dae1fd87d27ed1254803884de5049e1fa6ce734b894adb08b3ef5b619b18a298426dd6e17665413bbf8040346028a29c8e975d574396ae898985337716db8b87e52de80fc8102996f83652428917ff6ffb399e84b76c991dc892882e33bf34dfb0ed84912cee27a33995ab069bc9d4468944dde805d30934aa1dcbfe434716ea02faffeda9f0b7df083d0a738bd3a96b45a1c5bed586c19127ebe1abe752ed2aa6252c1afe271fe2313937aab2b98243915a170aad8e00fdfa52af16f6bebb2617bfadd09cdf06d07695a8cd0d76e1dfcccc86a83e9510a16d5a6f724262204c5c199d763d96ef9a134167179adf6e09af580fb2a76753ac0197ae096c53dcbd2b388c64c4cd7f5158d93472676766c59a8dee6ebcf6ca8b3744be790b51c4b199a8012ed76357e4fa5a4d869dcd66ff974af5efe252862c528bdf669ebf059edfd57c4923ac141a9cd1657406be03c73303366260723fa5edd76f57a467693b9d68c8cac60177a7a40b5e21006e3bbde28e0a18454a01758c7f0aa5f476e03e71589168047c5553560747711de041eb9f8720b3fcf302d63be4e6b7a7c863dab7e3cf3d70c3c6c0270bb723a795f53e0ab771713cb441d659825a347882acc9b713eee2b6e6d01ee3d7b0152196f4cf6d1550f1d6770f2766c60dda1ceaf5b2fe21f1da674451eb15b8b58544627d9f057fcc5285d163c1648b7dbc6889cb653836071bd4b2e580dfce825c5e68a58b6468db2324062e1d0ef55e578a8eface3da930fb2cf6bc3e7a5017af6e680a3887981fb851b3e943df4a0584f8e3bfd9be10f16c67c3773654ee8906bbb24c8cba6205b7d87cb234b1f4c253e08129aed111479122d9c3371c43db7a512c8addc516496a85e5583835f4710af40f57d8c6f7908056f99762a34ad838d37ef587cf22ddd821851e193563044c0d38a8f6b2902df7a502dea701e7509c1f59161b662d36cb94feb20700cee15ca5d8b0b5996e20e839e7e3bded536b17ae2b5ea8937a16781daf43dd25d41207151fc42352e5a36d162adaeb69bad5cd954dd02187fb610053dbd04231a6b50a640b7d6fced29709b0b6db45a2e200f5cceb6603d6eeb0068337d5d3dc0f782e12d9e76a074a62b52ae9a3dae80a30ba1cca441322306b7a066a0eb58b4f5662f219d65f3a08ba9ff7301a0b41c986c9ddfb05b3b3ee4154f5bad8def82f1e0794480bf56d6c02582034c8a2d9bc99536ad90fc9dc9f79a8d64c38367793410dbc25d52ff29cae0a51769d686eca8920fd1f9c8d5de9ab426b646c44c5b774dce69837b3bb35a58cadb3a43f1a49d6d5ff3e77f6b01590c42093c624aaae49d93eb601d2636f90d79d2a332e7b8c91f5a9d71017b1278c049403de6e44111da49c19180191dff216780b88c091e011f70682ae73ddc34b92e5379f9d886f01cbcdba858b4c7213289647723165a0719a4e67d12d68686aeae0708ce9afc1eebdd60c46b9e7fef25a8a80d422aa348a88f0ceb82498e04bffad5160d1136c5c8fc8b61cef003dc5e2c80b96b47c81a50315131dbf9990c45186636cc325649f1f4f7ed12d8c78f8e70e1d8afb35a730785a193ee04c67e55b33597632c348acf2d02018105bc2f7bddb3ab9defad388f3d2129fbf4c1d6a4decd361f170661016f3a5266d333541ca2940251e3086a6b6800df89749564b3c5f7b45230cf928da121e7ad347352881690302446ae3642a4de7e728bc3bc5bd52fb1b0f10f39f867e50b8c98554ef7fc03c2c205a8016adc87978255825d1ac67481384c4b06e51c51f8fa98a0c36fdf6b2810086372adf82665d9233b49b7cea6e2439a59c92a9e5b3d1dd9513fd496e73c96990119d0bf6821513b3340057ed491e7b79bdc73292db91d12eefb4e9feab56c6d97e0d01e3dc5c1812d88e1ccea9eba6b460d8e7fffeab1266fdac83921651b3decca35830688746cbd09112f4e326f9dd5175f0de6efd433555b64d0354be64cf192ecbc9d4bf0393b14348ac4d230390bb10c42d617ac650e9c8aed2df1681e919a2a18503de9b629c2271381b2f333b8a216dc189e4ff2a95886d66f1ba7b8f91c8bda8477f1ccb5300c485217197b7bfca06c6cc634904f9c4b706b62d98fd9d48b5850c7488479c1867d3a16869141bfafa5a5b4bcacc2dd1ae49cedb3e34ed9b5b364e3e143674999026c9ea396a78b928897e15f52a4da9f2f5288d1e0d87fe8b5686b9f50741683b47924b6b8a31b9d51c5229fa777700975a314396495cf1af574c49599829f5653a976f004e97f201d3fe0dc08baf1d66f3d77b4620d3c8315e751783b9f493a939d358a5dc4e0a7fb2e516aee0e9f9eb1e89d72492c59c5acfc1687aa943334fb4b545438ca741acae4e6674b37cd2aafe46f4418864e0d2b2e794082dd8b0c8109fcc53a578f098fc734d13794c9faf5696faae36ae2207f9fb7096cdffeb90ead0a309aead73888798f6927ef311b6d97a46ecc95053f7bdac1c087b47a0f96dfb6c87ccf50f30ec3f176ef2bfbb778c63b2bef650d8936561b0bdd9a7bb8d469f30984b0d83a026eaeee2c66cbb9950ffa19abc51f7656fdfc8ceefb5f048ab272b39dcd53148038a38dcfa56dc6664b20b1da9f6cf24c5c1c653b5f89a588d1ac7e3ff0a51001a3433dc2e6fc18dbdb68986db2cf53383ff206293e46d3669b1fe36b11f262ae87595b55b73d6405eb8d4ed47fd716cbfb78ad67bcedb53b78d015c40556ff5ff71b09ca08549a75a0345ccfc113841e6c9dbc717b5674833c3a98e7430e24da32f56d15c0cb0a334f7bcec649aefd38a5187673a9a6f45b7c76208d5acfd40e155ccdd0493592baeaa5f86782e0932a1a3719dbf2622cd44c528d813ba02f65f8baa452b0aedc873d3946ad673dcfc28bcd6ec3e4b20343f8c4218422c49b9ab3c02fb6e6f6a41a761b72a5a5677ce80262379bad22af24eca82de2f647e9c01c4b191838143d02b8eb91d27688a943b84a6e3a6753af07326c20dc1478f2badd45077d215de9ecb412279b1e0f227891c312e81ef4c97fc4487901be11145419a87b54c46a1d8b223fbbc14e2d63496e3128179e63d2b87ebb49c0d4e7b4f6beeb41c918ae4211928f6583a19643d124c381e69f32dfead7c0be82f5ae19f3190a1f8d40dbe60ceca99e9fb9e52528086790c357096a28e555c9e814efe76a8e33025d1c234c52be2193384e4a85f43f9103f4d112947cbe474677cd694fd38b13fa81e5aa7e73057236900d55f0c4dc198f1cfb17c81ebe94c326718503a2f0d92ccabc82baacac51879d246f5da24de41b55a8389f1a97dec8a86d6223cc806dd2e1bcba10b5e825314f3be029badf3e50049e833d67ee2f82ede029a4aba6107225435bcc542b1430834d1436e90ec99d914f361a621cca6835589700b967e62b387d12db2020734559166a4665bf29b495f8553831a3d0993ef9a74de5b02336cb7ef02d50be77af68145b9446df3472f776916dee44858ec4a93f165a030009cb22fec065e927e191b4c11ec4382dcdbf718b5ff4a456a69bbb77c7bc11fe1a496b739e06be873bd7415993a6f56bdc7c4ccdb9bf05a94d86ae72bfdad0477939c8727c97c4372817267cc8d308d5b6b2ee39a6f8b8a5ced8ef64d3736f003556cf505450f291570a0769840ac8265b674b1b8402c5d9729e940c1b5065c25a06303de6a98e0103d75ce6b9113144996572776baea1012c94f77bc02c0ad0b66df9b84e2afe066a79666123945e70f4bfc71c6693bef499f370c596059e6644da70c024faeb837f22cca4cd79732be51f44c524f73318fe5b58b1d5002025bb09d8b0dc6bf3dc74a65eebdb7f4e6eb11c2fc5c7f4e6aae121752d456b58da560dc73fa4e0ba64f4951636202ea53aaa4c638dc25a8c95ab8a21f3236e5f9b651e1287b1b775ca6a80f97723490dfa606937b0194b250e450149aa4f3bb961bd9ddfea2d43ec5983ea8907d5b96b09644e9e33669a6c3f5e2760379ac33949976915ebd25b42a0a9047a8a508079322f40ebf139ef2518c3e8249103792c38406a27bf350ac8f587fd4281961c23266d01d47b583971bc21dff0753fe61f577c38293a8946f7707ac469ac3e6600ae63e7c00e0aa61c5d5013a249e2d3aefc526409b605f86b2ab03bd221770d1196458b8c2683bb9a6189219628349c6aaf184b4131b8e6cdcaec4fb35be9a40ee76b7e184f85278eb69b594140589f360f5d46d87952d0928512a8f39f5cf66705c3347fae879a638a07cbe3da6c71fd51581e2c47ba17ebd2e709243392d1ce6080c91dccc1231d250ccfa44775078fa3886e624418904ec33e434129074065d3b300932425c8133e07b7952b25e92fc4a0e218492c9c7b2af86d4f8cb0f0cf73319a883c253d5899432cd53d8f45422ef202cb863b73247191b07d49c0a2f54354b723bfa2d1aa9ef1e5a7e61e6c0fb82ccf9e34fcf6e1fa9abc55a2dc5f914565b6e20eeb753dc6702bd580aa18013bcc44f6394773858729640b505593acad07f066c194f989362c64bbde6da9ffe6960fabced2d1168d38211969a857f5c26f4c29def3ac031182e7559209dcd14db355fb39a86ab92bcc7f18457ca43c4cffb69f2f6bc269dc09dd40205fa4fb9cbc677e4434b042217cf4fec31d70221e83ffeb0195191ac0c1cb95e908a0cfcc2a6c59be35538b3ead89eb873c4291d241bcd1d1c37bbb1a31a0ffec4be6304ce2dcfd3350905a84fbc4b89bc0aaf2498b4eb27bf92b6efa62bb6404f783a1948d92526a0adb79838a092371278ae6127fd00160cbc3cd90742245d2301520a7253dacbdc814b174cc45dc20b11cbc32448fc4b0778577b966c585fc2d442a0d94fd7c4bc93fe02e39cf52d0f5c2c74b13071af50d380335a0c0df2de60a870bb469b026ed803df0704d79471839b13b0692cb181ba92dd154c56d377aad809b608926a92a92d26db4b2e787c6d71df47123b7d9c37143e6b085ad9fd147a0177814021410b5ef0c13cb481650925c230c273cad81e1049c78297cc0a80d10f1398a5e7dd81e3d84ec3b29e2c6c9871fff71751aa5544c89be541adb5008d0413de11abbc2e290a991969ebe7272daf4664fbf53df9e74f26d925f381caa7d8d9829415aa085b66158f5f7304a0cb035c1b8059c26ab8e6cf78f24bd01a5ed33ff7747055bc8674c1f0ed7863d863b3b6132557b2f165bdd43e9f6cbae8bda6d6cf415491f383b48abeaf1f701639838ba92baa4db96c9340de14fff4bec2fb597f57afbd60347f6bb9f45eef4c0e99f0931de29556a8c8ce75d8d57cc7128917f61506975a9ebee1883b974d0f07533486b2ccd1e13887626a76a7f69a30083956273def434608c1916d5c227a536c527b10c9d0c746753f358c50ef559153fe51da7c394a47581ad17b1eacc06f95e62bf0f370a7cb7446aa6b4498b3d0690426a55a74012517b6843077088898854e042e2775c5eb6da339ab00657e79205a6f0d647b5ea7ab147f1bd680b37e27504e6fa213f7f4a4fc6211fdcc4eebe820d03e7e508a52575ccf1891d999d65f33bbfadc8c089539b0b266b4058f51aad4d982b267c27d5d3346fc2075ddcfa280752b1456e7b036fa5b917b1f17f07ae62c6b17fd22cc5c5d45e1dd204eb5e9c68af73ae6440a1e022eba2d1ee762f5c74dd9a83ed084a3aa4abad10e8f99be21da0e4bcd4aa24cea11ccdd1c245128091de51eb1f9055febf0f8894a0d82952d22efeb35a588a310e8b97e25e08cc41cec02f45d0d807ae45b80c6b3f353f0edbb79a489edbc3713ca011c8e75834570219ea410a89930ac9693bc4df70ae440c0eda82971b25ff34844798f2ffb82841033fbed47f4d8a580180a02c9ef204f4fe4419526af630aff0dea380c672aed4eb512d44af696618c3167b893cdf8663e9e201003e09e08ceba90dd3bbd2947d1e8d0797308112630c24a5396dc90d68dba816cb36dd930d6b527d787cc422819e40cf546cd8cd4ce688f77d19793885967e9c3b62a998fd691c4c5c1a2b6cf670e440fcf0fd36a56ff0f6488a925cb01d6fa661fd76ebadbfcdbab392230bf0a455c479572b74f4361850fd63fd9c7b3229d1b6615ec6c39a6c50af63d008c2786086b9788a675330f415b646de2859a5a11b1d375296221147a7d1d6f47c7aa61b43b61a6007c1a6bafc672bf1bd060f589dc8c6d0cf2891de0ace3a89a32c15587425a1a73ca1ffe6b90a51fb90b6c0a0bfb70e01f2c397ecf9352d8a9b4ae7a51f9aadf6d69c54c642b5918756fb44fe828778891f5ea5b2d6298c17af6d137f2c4230c96bc2650c040a729000ddee8d097346b9609b21fc81f664b11fc7cab7d9e6d56888a9d7415cb008c71d2c9c307ef74c3e88c52f2676170497f215797577b056e21e879ae21f9a466f647af365746d5da9104a7460423e8f549242e225e0cc05755db25968d5c968dc40788c9c0655f50a0c110cac690eb1f3a414244c17894005e2d1ff8f3cfb9e080cce53b4ca6d79113adf81d5120064666d1940b4ded5597a0f829582e407efaf079f7315d18c8577cdf6908bd376907917470c27d053dd533848b18f6497fa1c438b8f486e465f25f23fda2ff57f92157baea16d57d6194fae43d01f26b8caef9d11b4f65138226c3d5f8260edf1648ca82e60af4f83145d9fbb9b815539987f66ea433ac134606fcfbbaa7d2fc16958467a682bf36e1d729880af6f0301625d36971949bc964c54728542609a8180f277f8be971a11ca0c975b3d49c2b8326a9cf1365cfd939fd6fe5942bc9ba42e88c449d67fdfa02722373fd711ab43caec386cf8f64f239cc24de3ed85b896d2c3e35e35a2770ef648cafa00dc4528337f59a3050d76387af977109feaf23921c500a342f07587913f48b0ccd9e592e33f870f119a34b5011cc0739c0d323f2382e4f4687fd4a561059119b7cfd54ccd904a5d85e8cfa0a763c024d889f1ec84807331ed46e470e3cd82766524a43fffc41395199f3e788532a0d6499a2b2fd80bccb25955fef7d05c32fd7f5d4dfd1d03a353cc0c221cbfbc19b161be9523aa4c9b696d4c3090d6c83f103140da09a29f6343f95c7df927fc3ff98e32ca1061c9cf5b2b71421170ef8fed15097ae55cff63d5272a36ff59be0ae635ee5abc2cf1afabde708df20abf4b93aa66ff5583a2f4c2b258bc3832aa1da9b585442a7e7a1863ed9d91ff7783a0d82a0357c0ebcf72bf4429f98ed5a03a03b429a4a307b84822035b55913eeff303259b4098911ed8a79588eba2922950cbeeff9992661548a51f3f121aee303f44ab5da5d72e4722d076befddccc571aa9114a2e6ec0c426b5ee12c3b9ede8dfb879c6ce0ced9c9fa7d75d9d5a5dfb74e8f08eec199d2d63b140e9a1ca61449eef7472cc548ecbfa56f038a559793dcf1f6299b7192b8179d4b39c0f3a6290d5966e25f12195e0babfe27c550fc3abead9d7bdcbe42572179b8d7571b32e5bfacfcd983c24c962262b006b368ab426e8c41316f1703c20f0f3333a59f3b2e7adc515af6c7d0943a8b7e36bfc516e75bd3653a723f8bd6e93506b62efb3bd4191f4d4e557255f9c5900910304cba2e3762005d47e393ce6cca93743291801584ad5c44c234df4bc6304c9c05a5f25e0799fc7ee9510a4012e6b7961508790993b674eafb5ef508641b39dc91981ada69551ab4e99b747eaf33e047554ec8d08890114c6a123787a41228455c3f8d5ddcc81cecaee7814337370c26436862fd1fcb67d61b27c39da5a22c8eaa3946df767d93f5c2a7f271fc10dc389c2891c7aa9ad9b26b029cd4995906a8a2e09948ffee512569f4f7a7567dff3693ba809ad7c6b65b31227ffeb247feb5fa5776b302c9b5a2b0f0b2369e0ced87a95849a10bbd075dec78f031f3bfc61e52e85c64633e2d98fcbcaf46a8a808bd474d2ff844fcab695c4f30dd530bdbafc336e6e71ec454ffa46d450dd138ce9cdaafc3f4492f60083a2b39b92aeb452cede7ee34376ee49522272180c4bbeec208dc3e23363328d0be9f6cb219455784fca3aa79b9c4a11cc84ba08ecef032c9cee34804f8f9031c247e23bd60c362484b90b22682c328d7efbfb6489db36e5fe8f3a8a2e65bb22415606f3f0507c7953509846f5d4cc4ac52d1b320d791541542e1a0611224b5fbb4e5f812047adb6609d2f0a933dfb1a44894f8efcd8a73bb1bf2dcd1f2554b92ff587077023fe5152b8a6d3f542fa55f9ecded7c785e968de0ac10e92ebd5d0ccc76dcc1cbb2d8cf0c7b9891e65d0594cca8074bde24efdca6a1ae6f5e738ddf78c57087ac30540ee745a10bc50439e5654487cd1dda7739640456d0fca1b2cf5371fb8a05f628115de0ac8b3fbbfc6295c7a9d15caf91804766e7cb3ab2598f4027940b1199e17667f6b171698e76231ee4f379210a61c15a195e5bf958f6ce6d06845bf725c854e7f65f1132463676618cd3d671dedb0c454db2f17392f77546206a016a9ba3239ee98c9085b2504df3103454cc1d7d8adc86d687bf9bed0b22163c599b3a97ce5d5397739734aad2a3ea59268c6092647a6b597b41265bd7e8c3812dd0e20b3318da3e0cfc86392d2bbd32f86642407b932a9831184501806a79f3e5ba903f5b9616e515d8a481cf002b2b80ca61ad25ce5f6e31fd2f98f85d40d665b499f0ab5b8447e491ef047a011cc3ca49449b435c7eb170f380342065430934530515a88ca6a7e26a0100d8dd4af6c69176ad2c43cb4094923fee5c0c06f356820925d4277c8aed69e4746292227034896864ab586895ee376004e264b71105df14622daeffb2951f4298d2a99b61d4a5237a2878b7b05060f4071455b2986805822052ce163b6aafd8e944c62f4174f3847d7c4911e1b6343c91a06462e05e02cc32a0a519ba99f8dcb7dcad2630ad7d6a75857629c56adcdc218212589a67712bec8608242acc154f0c9ef76e63b1b975e4c23f49e4f86ae9853be20db68b453eb32931d4ff500f2b099667ddeffffbf4ccd020f51b26725a1d87a735e9794436b446d51be75b5d98c707b1376aebad8d1f12ac3b842e81362afbb075af11f5271e254de0d13dd4bc538af2a5f15047ed62269184abd61129a464faf245917c491fd6f343fb19a6a4e1dc4c87f71d9bf81275568a2376b7c2bd12b2e6a4cc5776add167a2c6156ac02b24d0d7952e41b180a14ed43b49e40aa4de12bd32725027e10c5315983bcc36f7a777db224f57da964b959969b6f34eec76e962a08141a0251b05ba7a14b9a252bb8e9cbc603338bab442e5c9efc9025a79d22482bd3b0f832ebc27648f58636e3d2bad63c1b9f399e90d9c82d4a1be5cf55bbd8ad0718cac5ad70565aa5dd623f9a09038ff7bb748f6e9a4e76aa969b92dcdf5d6d422e254a30562370cb86c36fd2662441681734a5136db2ce486ed7d2e5df55f403b46ccddcf85d023dd9f5642b56dba9bc406078f9a77dbbecd6d1da4d4534da6dbcc50e754e06fae8efb584c1ca302484532c8b6ffcba8365a80b05bcf5e37efe9f7b18a7e3c89e5d4d31d81a75722eded4cf94e57d41c6825f7433b414ab599d93bf1efda78fe5bdf431c6340ec8ff46f1be76a23d25bd3238706ac1db6116483332bec7b5c68597a8543b50754a8be30a2190dd80d4ecaf821bfce9745e3e994f84a5ef28a791597fe0354eacc0b93c0cd003671de34f2b4aa5d709d2552cc4cfdeeb9ba55e8cb451a4aade229ea03809bbe754ca56b51865582c7b16fc55b51eed9143ec1ff44a395010fe19ed4b0634856403908b5f29883c4f84cec33af1c776335f5b2d27df7045a01ee833519d8ecb27dc7c356d6a311f92f06614cb25960ef6a74ab7ccebc2202c88b530a00a6db036c33b44d75ca47e697ac73cba8d8691da6083a0551984ff73c3456a6a54cc54b280d99c3069ae0ce3f02df6b25c4f6298920ae3262c69589c89f19acae4f57d9966a560082021091ba55162eab845bea4d421dc15ab2e4a48272b4a3a402190fa758e49aa9c9ad56c19b94ed8b66cadc26e79a281d1951d943af73837d599c55862091e459c9b8722c96c13b32637dd6729a422d5725dc75866c0a1773e249876b3cc2a867645b8325d67fcb4716e3422c93bf4e56cb2ca692d44866eb2b749e15070d91803747c80c6dfde7705ca6f60087898ca6e84d7771396ca850b01ddd3c7ed2841cb95e295e0dad6bf1ad07f740868c9792191d5364ecccbaa497517ceda3eda2d6e3098f469988bacb6498e0a3a0d180ba63c385f30098766a18d5c208c67e7bb5151cb81c880d6cab5b56bc382c03984a849a6b1080683136e829886e1e4da235fca9c69ea6705f15e253aabae1d5713569ede6219031effb5104e98bc54024e5803f316f6f8f7c7f4b9506ca9614925d532c0fada5c8aa1a6cb98a609aaa8dc75c539790a9688a06deb15d42781ce0e19ef86071a5422bd716ac4621971b9d18fe0b029709d203369a8b2cf91793fd0e5c874e2054516493a2f5aaa9b08feec28a99e9a86f70ee814bf64dc0d02c0c23e7b6117f56ccdefd72e846fa8194c697758eb2e39c0007651b0910e286f98866d006a7f0f1daa037b8370d0600ba4b5dbcc3a3ee25ca3ff65037ae9d823c71483c67dbadc687e6135735913db2e2cb2697efc8429959947b11c227976fe6ea4ef17b4cb6882ce49d5385acf1a7444bbe4048f5d8a97d2fcab42987048541e183bacaadd9d82b01bbbdf2379891ae6ad6414d81df34029ace237aba81cc873c9adbdb3f698899b7875751f111984c679d1be6baa0bc79f0401eaadb1d13da3cebf7da05362502b150d9525c2061381d6bf024b91487b616cfd27734f0bfe58bee3ad578882e70e0036aa1699a49a9cfd1d6768d548cf771236c3925c9840fbf960eedcb19346ebf9aa97c47b9f88e74590026e5fa0a492835f358a8bc0611d9b9130ab8ecd99059a4d5eb35a18e9be0785e316050c3480c9efb480b21c530b01e94fcbdb1704ac0f2a4feb547a32048b9c5a3dd405aebad03d9f13004a853d8cadfaf12fdd84c636b7f237754f5a4899e93fe4b531b9e0cbb6edb4c25fea316ea729cd710f049fc1aff1d3348ec0c30c53835cc49b2a022d9e3153b4d5c0a2bab84e17b40fcc2384b7cee7283c332f5e751b1162c1f8f5aecaa80fb8b0999785ac49c9096fcdb264884e8e00afa799b23bd69fb3800cc5558c33f2aa88218a9197cf5feb9ee3b27a64c5e32b5dde67955e8497e3b429dfef1f4c29990feecf9b00f0f32f818cf789f89d03f49c90a12246bc895531fac453ed92f4d4df1c1a27d829a574b3827d12385b4ed4da1e5e537494e9a929ba58858ab602e6cb36b5d82ea2756c2c204a605cfafeabd61c729a9487a70b05b63d2a55883ad4b7f62f67ab29b85e7a5ed25605614ebccfd423eff83b1386102990feda815c0e5fdc9c44e440948e93d0d42519f0dba3b62430f2c5a7d595a3e09f2e0388dff86515ec45bb10593990e769e7731dcf203a82559ce526fb9478f7afa201ec6b3abe946f4453aa0c3447b1d0d512bc0739b2959b2e7e58c67dcae6a84da2c8ccafc9538a4691f33ceec74f4992ef451a5a66d11315162fa6378d796ccd498f44454fed63c9d7bb7402c76eea5728330ca929ab87a622114b205f8b6ff871e18888ab95edb4c5078393c5f6faf34ddaed97f445c142c96604bcca4e100f9ad7f79e96e3c4ae17f4f7caf8b1c28c152ffe520c36bf8073c4ecfe5057b9af45dc37fcfddc633e9b29eaff7dd2ed16783555d2e07c718eb418b805d631ad2393dc06dc385481b2554c27001f14a13886a3aefb430ca0ff0ae88a8050773c04b57a1498d066f8e067ccba6db31f43ea450cd05b5b5a5ad1202e77c006e6b399b7fd09bc7f5019965f4e7de2f86abf023301aea538046689a3a2e3f7c862fc364f96fe704a70ecf267ee7367bc66ac3b06e9079e269c2586028817c4ddf092e11a2f0400dd3e08a8588f24b1865ee2eddeac65793d6dfef5157f4d934650fc938c6f77ca440d689b6c76f23544f89ba7562439de0991c2bc98d218209ff06d40f7e02bf8af6b60259b6f2da43c0349b518c2847f0954f800a009964549795e0feaa5b219073ffa4045ec1c1973fdba8f4abdaa07af742ed4d9057ddabdfe07d1d6d5820f519b5c33c7271f71699a90459337bafc610e259d2c41b6b88610ec390fe69976e905eb53d6585af86b7a09abe453d87fca735d6701d84d129a1735d57b94104759eefe094773d8c2aa3b6355c8f2abfdd88870eb030b4ccfed7e60caade345c073baeb7d8ff6244cab6aab68b1b23c22569ea109273511d3603549532733b4a29c5f3f3b9d2c74cbe1e24d78a38aa499d6dec331e2853737bc0469221da2caad2a993e66358db514eb0b464ace04db7836534d79da5b083ce323a03f0ac08772ca7150709f5c0f0781b90e0635ee4b3e10a9c97b3e56a697a7ad60b46fd843ef9c47c42838de063b485828a746d23feb5fe9ced53246f5c68954e6d61d7c0565b0326d9f5a31d892031fe838eb0951403862956409e24a5d40c7d5217ef4ecabf4c44ae33e2685e03ae70aa29da511df4ea2e45118b0cfb2e2b7d423a2cbb313c1daa5c7901aabd9db1e1939d2fb61c65e7c923436c8193401afe4d114ed481ce308e4ce342830396fee37dc8c8ea876b3a09afb64936415771c5658a2e965f650079efb4d1831f70ebad7ffdf76972dace238d9c527507c10253c55ade027ab8af3a19060eba34880c44a0131586f6b89fc9a269d08e4ed4debf500d39e2da63784ef58d0c3130c55e1001befc3d1bacf503de5d9d6ea5dc0ecf0a776770c45e3ecd515abb16702b8024512ded6d7852cada0a4ae56311bdfc2469abfe624ad337eb113c8b72054805ff5aeb8fc37afeedf6236a641e8ec65cc6607529e5df2f357502e7515a0693d062fac077eb05e5583f8a042b4d919b58520d7bdfbe8c041c3d61d395ca21c5801765797b5cd277e7e3e6f6a3667bfd54b3188645c4b32fd224f6533c3bb2e849522ee224cad226fc54819040da2e558f78a1336118d83baf025ba0fcfee0b90d198a05edf2bb235d1bbf2ab88a73140b841ea6c8591cf9bdecacfb4c48c267b03a0a58521c8048f5f365fe353a6a71ef8c85cc331d469eac7e93500126137f960f9baa00d3ab3d99be6ca03fa3a6bb5fd1e1a32a43e9982d8a58d39bd0364154125abc1f252b98bf5a5fb0b170d3c3702ed9c7a0f96bf9e39534359f85257f2ff249305603f16fcc24e66dd441e36cc547bb68b05dc31e5ad0cfb78194943d30d0c3866ee448080a750961967485911259eb3fe8c94adfc7a27ee3ba7bd92689c8fe1e8cb01fe7173d99380d83aee9e2b9647c4e5a7ac76aa3d402ae0d1865025017ffd57880cb3d602a3b02fcb0caafc8dc2c60ebeeb73eb1370cfd5bce4e74330c0c2f2b6eef45963ba1cda096581db0da60764fb61febe5d53fc54010b41bcd2604d2ddba53d6ab79c2fce3e79583426590d78bc512a20cf3ba6d0ed852e5626e8f99c0206d429eefe6a5907f768e0f644fe46ff7e3ddfdcec384a629e1ecc310ccefe22239a56db565e3162200c23a7e1181371e9c42996ce2de53c58458599d171fdb50960e3021e495c91ba619ee5330027dbed107dbf1b6ff7b2f7dbbe74a1e5ab56af39da177452ae16bb966f9ea9c075286647ab4bc37b8c201fda72b3bf4d1d2b6b7f57c3dc95fe5b62383bdf835cfcd541ba49f7d7f3413a81860787bb11a8676949d217cc58a7c6f56895ded636e3931dd35b538e494b58678ffd4292a0b14e19c4c9584ee73dfb9fbf1ebbaa8441b3637d11d4caa316686ea36a9ea9d4117aace27f95acb7e176dd4ba9f6d934c479142fb8c16e7a7c29120f920bca136116b783d31c107932cb784d37f09c13bed947ae4dea7706072cf2f40dd782ed099361e85fad0629f4dfb3b7fcae39719f29755db918c4b76f378e0602593152782ef7b6e09d2ea07d3eab79bad9994f6b3c7c9a6382ec80bce1c089c3eae8b66f6e7b634a6dd60255d38df1af82eeb5a61e37b7d61c4abb065019a311aa6e589e8bb70fefa6083a66ee0d30b9b0fc55fa0bcdfd499e5c37bda3aca12511fb747f836c6afd7404b68fe4fc5e7a51feec40a89f35508dd8ec8f10d22b8ff874de5577699cf5e287b00360987fc7c95997288895417e2fe259852d4db215f6962b7e93039cbaeb598873ac0dbbfaf468217213db3b8537aad4874268652837038a74f05f518e8fc4720b12c3169b2e4f0ce398a485ceabd435ce109a3096b79a0a5e534b0b18b4457e3c0f04f829cb2190901b0036512dc7fdd27a8b45d453c40a1a28b26f46abc04aa17fb47b8dbf52a74b8db1c9bdab2cc4472b975ab46632f881e76a208fa7c30a46f626c25b4fccda548254f9538c7037bf837e68cf467d0802f0659956a197d5cfc6035dd159a1062f1f2b606b9d21dbbff8353cca54cad73f9f20719892c6e6f49eac2e7ac2c7c4d3620393dcf4d7db831fc94e5307c4ad5ba03688ed2ae2191aef1dd38e09dfb84a79b73e6c7a39950075c9fefb71e6e18c700552c4345183d0ea0d227c32bf90c6c9fcd5ff5c63b0f497e8e26c03bd26690b99668656d1c08b923bf95b1a9760c2dbb845aa57641ada383c128f807ae1a19656f98afd6da6d5c03b67ef7fadb40902ba79ae8ad40957e41bc9a0c964995c96c9aa7ee9ad09356ea4cf0f327363bd61d9edc1bee40c3d7b797d44a796a5d45cc7a45add759f9dec33e7c7136cc761df1848a7eb264551e0016bcc4aeb96fe37c64d2ea1be3865e75c4032fee1f554bd128ed832d983de7d7d54e58252dec762224092dde57c08232a61d9fa172aef9be5c7a282f72bf481e44da92e7ee18969ff7d7a770299795704feb238decd53e34f72fe1db61424d8d26567f2004cf7970cc075f9f1212449ee0a1f57a19aa0478e2b9446114ffcd0c3c49036214a60927fac1e45dbed7ddaffee046bf7d7566df98cfebec14497e9dbfdae00193b97255ac28ec425e908a5c969325dc21e91527f60d0a95499c95e6115b3b7fb81f88120a51fbdd6b2d6c6ab6218cf43c73487d4866f7260c778b3570b086b401d5ea852d51e5601d014eb14fd7b87e3add6db645f45e123b8a77c2b6e91cd7690fcbd9a77e64c236dc74ff23b2a4eb49d5a1d9a6b92801f191b0fc055882cbf01fce355bf1850f87018aaddbbb5a27e7dc3fe9f52b9951f360f2fba90d1508ce33987c729cb3028991d9e780687d8b06e9e3149626b5e957466a0fddebf21f71871cab2cccb4cb6df068e1328a16fbe119f262d73943f1d0bd6f93d7e1a03ad0fba0ec719e7e30f909ea1518404d6689e9a08e3aef56f0baa5812728094a1971e4ff57b809a9cc25b0052af506fce69e563f1821d16aa20dc2fe53c25973b1341831671ecb1f480b4fcbe6dab5d3686393377d5d8651d02df0c0a61df373a0778147c1f0dad3372dc0b61f9a1882f74f56dd861249ec011d8ae668830ffa9f71280618d43a468433e9dda9ca3c61843771cd5f72fa1c4a84dfc8890ed1d2942f6eb594d88c2a67978f10f050eb905efae38bcaaa5430c796584c664a4a98d6104fe6dbc853a2f67085c3a5bb917a155ac129937df24e197ea8caac5284e45d4c3435f3c3a5904f0fe264bf4f8d9e2827f04a92b8a8ca828b01d59ebf8c4d12f64af564ea53a9bd93c273118c66a6b7ce4bc145b46df232d1daea41f8ae96701adb148618d9b137eb8b6b32af6abbd593dec821af5ffc6a14fab893556d75260af9ba48e65173f32bab22db4e3790032d7fd249083338bace8ab1bd82c53ec211a3df7bf239b9f602b83ff26e1f2ef0859bdcddf9f3432675751546d5c8d06dd110bc8d63e7c478cfc7d63039e443ccc5fe283f6c60ecfac4bcf61c3e1ca8c837d5f33cece6def60c662d015665d4ff9ca9bdabe55280c721c2fe27e6deffd9387662b00c9a51b7916692d221cb81d29204fda7744cac65b05e911445158061182d123f573f897fd7e48bab6b281e1c8f397e072a573d62cb143dceeab4dc2cef3f1acd50218f72d06dbdc3cdd2186fcf9c753f905f5a6a382fa70d1aa5a59b631b1bfaae7f48a40dc624126c50792129b47fc63ea271deb7f48a1c8e975ab81ce9f3cfca585b63d3a8ae7e46e860aad2aed5664d12df8838d5f1e17154be7e7b8c99d351a061795741024bbea3c506a2c806689418a700447799dc1968d48d8624116342043e3872187628f1349939f5c24cf17c1d4c9dc0af002450aa5a5951bd486c4ebfb90c7aba880e2d1e542bacd9802894d5b2ea4e37c9c5008c83b60ebebb39e294baa3ab87a0bacdc1ebfb98a72b26331ccb69f467689e3d9be5df836c55ca1dc02fab0b54483e62f0b54a98d0176ba794e859975741eebd2cef586371608a7e447a5816fb18e58a69476174b985b5e1a46331be7677d94bb1d3c3f0be201db1f68b7891f50dde37c455d2b4a6464df49f33a027d46ccb1841e5d949e6a45a37c185dc88057d32d4d970f01208a8f6b9148e6d8c054177439653780ade95d4b172e3d63eb03797d0b59a1e77873eee28bec93c1b446b0020309133909f8649d46ca443190733a1389aed61ce8e3f3defcc847ad656b15f051c9966eb04ec8294e61863425dd67f934bcd1f4d73707608eed8691c83c1da29a68d282625c571de2b3e7cac472523de0d93f72af877824dd9ac3b2cf043e6a43c7b4bebe26fc96d695b402018047713ec5691f3c2947a5e13fabbce090794e0557fc267a8453e39d4bca4241609d3b87e27afd399e2318f7b21a70ea1fc4b4f652ddd5ea3cb3a621dc9e88ec6fbc30575909b43fbbb75df06c67be8e545e8caad30d1fcc576acb6941cc2ca08d0255f30788e754d7f486b4f5adc1d2e99a56bfad1038b10ba9eed3173a7f5b67ea5111844893bbc056aed3d024f47693fa8082a6fd42b7889580936a6830c1cc141bc103999249422ec786deb4ee02c2dc78171956da786e82bcd59b83a2039c38c2e5802ff823e31bcd32e0375f3cd7526de586c52698d37e60399d357a4920dae9194fec4c66e19c259df5a2d3e0dd1a103917fea0a2c71560cdae449fc90e12632de6d1c642d4f2d8dc85b32a78d9bd36eec20fd67c0030053ef1dc7ef85713e3c181fc463e97ddd27019fcc387cb7a1097e1111ff7564f20738a0fa25b489bf430efe02c7da1035a78913109c4071bc2644b641fc0643f305154de1f86a13347346d2f7742ddcf2bcf7cd36a3780a1730a03cd0da21aa20a3987c0bb784a9db2dfd7374b4482e1d29111b3121e0cee68c99748c6bb62c32aadce5b540ae453e3e098df888184c192865fc34110ff1eec590e80d8b841e5a124de23c44926978b83a69ff3435927b16c101aeb095251e7ffdefd2b2e417d666b33be6e40e3a25f4b9b932397a486e0220a0bbe65b868e28e0df0ce2b9ad6917e336f0c56b12b822c74bf2e64076bdb19ff49e5090394c9234621512a8348866b0a1dd274d0afb465bb8fac8d7d4951190caa5f7b2efe6f3a2f30df89b9a33f2140dde476d2448191da1d135e2b491699630e72a9fc2166f718ac9a6e607e27fe98e836533d168f2e47695fd08883bba9c536abd38cb0409a55950e1962069b0a0ffedf735dc0ebd7d20b2019a9bb99d325643856b0fa3c5472a3710b202e6a6ca04e1277c4cdb2f08fb28bf3db7f1fae32c4664c6a559a346246c18dd9595b2e2c4467281ec962e6665bf97db482bc28b9eb07868e32ec57fa6e9071b85339cfa1891cd1c3c6d0f8d49803cf3de08aa326e66106fae629b628d54bcecb706b59284aaa565e26070865f2495182903622de0820636720b50c61261f0e3daf28cf6628f3a814cd63eb11ee5a3febcbb6d67f571149e9229dd0958b648f091aac40ec65aaae1b323102d94e186479d86de0e6bd990500e400ead65bc30b263d4e20e51f43779ebc51d421d4482e124d6b53e90bff2e70189b10c9c333357b456c114c014c639b080a79ae0df87745e52a794d38f1549e9f923f910a69bb4d6ed0f621150010c78be831d2c0b2fbe130c6220e9333889ef3b39805d13464b0ba3ea9e480e7450ea0e56686ff8c1a9eb405425d2fc635a8143b8cfa123b73c694c4c1d93d662ef6bd362651cbd650e16225e2f4bc44c258ea9053fc5eaaf5acb542c3f83c4d8e47477e3efdd6562d403bf5345a3b55dd17423307c18ef69ab4bc846e9cca7a51254765fdaf94ae42febd3875a69f2a5ba217e88781c0397089c3367bf1b02223af5284b27f8f57b132a944453e1dbcfce007a68623bbb4e43b79b9a73010dc6fa12678c0058ea1908849ea222941426726732419f3ab91b3c5b408fe7f43629ca360927a7df1bf49c1c1eccc1f30bcc839a86d7e54edca375be862ae1057da12571807e28a118231beb87cfdc8924157f002965208af901a81ce224d7f7bf907b202c5d25b046a4138a72d73a113bfd5af4fbaf226cece8b0a2e9fb7c92764dfeafd41952f283709c2e8a137ba162bdfac3ce88c95b55a2e9c91b84b33df2e437e8082beceeafa3e0745c9e8f714706fd70cb703a945839058e865e99bcc4e666034fafe4d2a86221900eb117f55e40e8e64231330edb62693c63fb95d81a4e6c038b0ccebbfc17d657a168cdd1e9217f460b99a96ce4c2149248decf33201aae98f5b84eaa74f0a8b89dd8953a9a79c12597fcce897ecba29ac79325ec2d12c0534da7a6aeab549265edc354c0837c580c3903f9f99dffa0258c6609fd22a6e69cc044b5f64b0d25a6ade4074393c4875b93a2a16b8638755615c7ba47b6b15a7a3c6b6b499a4d1106e14f079d1423f0dec1e88f9d1f3969b0fc7dcd704c405e071b5064900311cf6b7ba503f46d5df9ccfcd1ffbb5387388dd236f4f9b0379aca1baa4ccca1de8bc232865137e69d28862f91a605c91c911981b4a7141a115b79919a0bc08db928a4ca63f9c4d7225b399a05805d099c4c8a1aa2a069529b9db04834910f9afe9b26b67732472685efe686e63eb8f674a7b8706217c50b9bc27c6c83bfbf5d938c167bab7247f7e692843f3f0c07e098917f9468509f3d8e277c59860a58b1aef288bd9cf2a85c088f9424c0e39d6acf01a0f1e22d91b053526543fc45411f267b93343d26a79616a569cf932215468704315ad1fa8a552afd5907a2e1e6ca80b4f7c589d4f466016d1e8f798f68b92d6a1777173b49c4eaa4a44a48984648c1ffa692411b7f86e0b170aa6720a20d840391d9eaa2e1a9e98712469b4f782e2e1897371892a54f24e2a4b2b4ddd38eafa1ebbf3012f77f08d958d300e038b9a266c43eb85c7bfa06ab7e3ecb509d8ee64d1893bea13ed5a4412d8b9a5f8ffe49f9dacdcae2ec62f0bfccb5f2cf53a79ad586b0606a5c76d3fb7ee7841abb198cc22d939db930d40f66201d42baabb0909f0c812c7bed933bb9ac0d9c3634f3350bde8199ae549a67acbabc49374ef3736fc8dd8bbbe46b4e794e34a1a5d24d150f44a49e6a1f90534a0c9f08343395128d63f7bb57e286a7beb691dc4bfb545301e9d9a50bf864337dd7b225cdee8062420c3b4c7bf80d2faefd46097059b7bdfcb3c9658d71ac4e42ec4a031261f9cfe368d9defd56754b04f5418145de65c1ea84467eeff5f2d7f1132a6aee5e0788d4d1db723f6aa6b428e015b05a5ba9ad2c80e894a0b4fc80f509337905901f33082806122109554fc7700ac34128468d9d9860325eac1219ed811ab7440be24fecc678a91b8475a70756c13df1e7ff04ff260e2b9881ca633d2291e39e204114eea3ab02a845737f3c0dcc71573a0bdcf5a9e3571f7466ad7a1013e18c01e38fdde8084c2282d8131c8e27ac5d5d281f876cc08a5e90fe487d41181a2319d74947271e986b793d578f311d79fe88fe0c60331022261e53b679b3806946a7632e0007ba2fc96066b5d9177f4921c78326edeee1a9132fee1817ba97dd298b8759fa7b6834d4ff463087efdcc29c53e304a12dfd5a57d98c49c2ccb0431794143b2b7f0c718ebd4d98760d3550655a38237d52ab138655cec5c4ba187359cd7c29d83b0011e45dcb659a99dea8be0e9e9d35e8b9eef0cad8eefe3400e10e716676e31b6d30992ecc6f85f774fba7a2a24a2bae0320f1117a2815ea1715bb34604a2c503be13dd215de35c47d4c4d41c1fc5b661e6f3a60b33bf8158b697aa0a8f11cf3c0f9c1e3f789a404fcdf59d4b8edf1f0d96013de8a51149c3f3c2bbd1d4da6397ec7abcd02dd878cbee907016d6b99cab7f2eb2682366ebe8def0c9b9ffd28682ac8b3f25b3dff231e6c5e96a2ffd0112dc5b6a5fde1d2423ac8e309514f71343212586344b143557b6cb9f28dc150ce880c6db8ed830f21a5ca7b77e4c79669bed64bbc7b1240fe2f1d2754235430b9c57f7d7873b1a6128ac4ba8f4286ad7bade497959e57b094c0306b9f3af1077bffa974a82b4ccec032dbe4640ac4dd526b4b66c4415dffd975cf79c0792a124664eb6575539676c5eaba5b918ddb65605de7c5f01a4bf620c7622436c3299d3d5afe66ab92e67847ce07457dd6e130a10463c457ffd67e8563dd27d8ab3b97380a1b2fdbe1f33ffe24307ffba9989ddc2fe053bf477694af974c9b606d4b6e5b2798020c160edbf4976d26ac020670885e575f99b28b3ccb61b04a387f92e219b39d679115bfa1acb700e77151cbff9c6d9c2883439fcab36bc13776472729ba231195822b8a87864286977e3bc076259b837653af945d03f76ccda6dbffe92c4595db461e6bfa6fecb18bce2bcf1c6b543af30c6e4d9c76d5023949ad273158ecc22c7619ef83f21a6b95b9ffc68d0ea60471c6461fb10399ce9d311f13e5df8bdabe0f'
	}
	// Its Shake128f Context
	c := new_context(.shake_128f)

	skb := hex.decode(item.sk)!
	assert skb.len == 4 * c.prm.n

	pkb := hex.decode(item.pk)!
	assert pkb.len == 2 * c.prm.n
	pk := new_pubkey(c, pkb)!

	msg := hex.decode(item.message)!
	cx := hex.decode(item.context)!
	signature := hex.decode(item.signature)!

	seckey := slh_keygen_from_bytes(c, skb)!
	secpk := seckey.pubkey()
	assert secpk.equal(pk)
	assert secpk.bytes() == pkb
	assert seckey.bytes() == skb

	// deterministic testing
	sig := slh_sign_deterministic(msg, cx, seckey)!
	assert sig.bytes().len == signature.len
	assert sig.bytes() == signature // PASS

	// verified := slh_verify(msg []u8, sig &SLHSignature, cx []u8, pk &PubKey) !bool
	verified := slh_verify_sig(msg, sig, cx, pk)!
	assert verified == true

	// the facing public api slh_verify(msg []u8, sig []u8, cx []u8, pk &PubKey) !bool
	verified2 := slh_verify(msg, sig.bytes(), cx, pk)!
	assert verified2 == true
}
