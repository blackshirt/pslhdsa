module pslhdsa

import encoding.hex

// shake256_128f
// 71175c346898606073adc3c823742789a47f37a5d2cf066522be4f3dfcbc141044421141a7d1841cf92d787816b7d6c77d48e8f30587e04ff4050e7817f4830aaed14f80d5dacf63e81d9fdcbdbc48d27cb973222164bb46dd24fa468aeb8400c987a1712467be1c0197ae4ff94da5566c1bfc1c88675b2df323c773138b7e9352505293e1db544bb4c2405196d1aa82ac68db1ecb07b29124ced822080d215924389e5e8ec8b149cb441309546cf15f42833f3d586fded0674065744baaa9c1e6d0be228172ead974bc639faa6cc0298402287b027c579224702eb031d8ba98db4cbad6400a216aeeae2e4606c855b4e0891a3a4d18dafc7b7a4d65323cc4ac784b18013fef0c425f812d800b7b8bd5486144e02379ae0bad28151bed3ce2ed0b5512100a2615590906abcf406cadef668d6ca17c2826c19ddfd841ba960f2ed1011fa1d97aef566edfde9f6ae78f9707b5a84eff321a59ea6ffe06fc1f9ec1789c5ea31a1a400416623f5535ec7d409440231b4bbf5ce88980b0330bfe5b3963d502b453fd2ee9197d5124b2b803e8a702600339463ff94a91bcab26a2ee85dbcfd0acdd534a70d4dcb2912c21bf7295f22edc102e320fba36acd3350e05b2eaf063b5a005fb44cf4b0333a2df2530f9d886b2ade35b1c1b528f74bbd463ec5099308b95f3829bad398fd7aed0725620fc4a435bf956d89713a895b39c5a585cbcb63ad23761fdb46723620daf32cf95f149cc88f04383410dcce8f0571d23a1d3902d3364467829ee37f3e2d9b520
fn test_wots_sign_sha2_128f() ! {
	c := new_context(.sha2_128f)

	m := 'YTwkwhkyJG3PMpDWlEvRuN0BppYASt3J'.bytes()
	message := m[..c.prm.n]
	mut pk_seed := []u8{len: c.prm.n}

	for i := 0; i < c.prm.n; i++ {
		pk_seed[i] = u8(i)
	}
	sk_seed := []u8{len: c.prm.n}
	// SKseed := make([]byte, params.N)
	adr := Address{}
	// var adr address.ADRS

	signature := wots_sign(c, message, sk_seed, pk_seed, adr)!
	// SignatureAsString := hex.EncodeToString(signature)
	expected := hex.decode('5d6b15ca78bdd156fbb972c2207016e1c829d861558fbc1daab4f3eaa7eac28e89b9248f6ace1025d8dbebd436672ee7cd354903450675ceffbc6be1fca0a58232543ca4b81c6e75c87b26d97e1752468b7454de2df0468818fb379ce91a44517402c3824450e7e10b00675a38bff69202640fa4a7b31af12bb4bc995f532c722bef7b4fe4cb814047a07ccbaec93fdd02bec3f9940ff6930e6d629a5af971685189c0d89ec78cfcb8ea439905bc466a0a2ee3788a8916f6647c0ef3f70d835ef7f5daf2c50a739ef03ee7f582a7dae4628e0fc1c9e037a34ac864b665246afedc70c79a1af132f29c9d15a322e43596d2011d34e267ae7ca853e6dafa25717b251f035ac80a74b614ff748c1791c8c360118f7616cadaf7d590de0aff01dac70d7e72b5e7a47126c8b3d524eb711a8c1964350027a8081ee99a89de7ca7a5d16360936eab5210c1672b53fd52cea6fc6286a7cb75105d56a744cf903902004ff413146132768b5f004c7264b1d69cf6fe3d5fe4ce9e7c18931bec44f714a7028bbbdaafe3b74b72ab82cac084c8a7020a947a540eca3f4e2de3d6640b249aeafc178a3e7726bf13b4934d26e08d12fe017f2f75ab010da1fba6abd2266297585d342d9d99da7eb8465535072647e237e2cb69532352cfa6b1ac442d57e408f14c38f5a94cdc46b5efc88785348846e754652f13b214a17a41a7c5fca0e61dcbc24101fea1b393cfe055e74215b0f043a1620dbfeeaf88d7d0a5f6b797e9bffaac949b574bcec9552bfbcc9b1a377299')!

	assert expected == signature
}

// sha2_128f
// 5d6b15ca78bdd156fbb972c2207016e1c829d861558fbc1daab4f3eaa7eac28e89b9248f6ace1025d8dbebd436672ee7cd354903450675ceffbc6be1fca0a58232543ca4b81c6e75c87b26d97e1752468b7454de2df0468818fb379ce91a44517402c3824450e7e10b00675a38bff69202640fa4a7b31af12bb4bc995f532c722bef7b4fe4cb814047a07ccbaec93fdd02bec3f9940ff6930e6d629a5af971685189c0d89ec78cfcb8ea439905bc466a0a2ee3788a8916f6647c0ef3f70d835ef7f5daf2c50a739ef03ee7f582a7dae4628e0fc1c9e037a34ac864b665246afedc70c79a1af132f29c9d15a322e43596d2011d34e267ae7ca853e6dafa25717b251f035ac80a74b614ff748c1791c8c360118f7616cadaf7d590de0aff01dac70d7e72b5e7a47126c8b3d524eb711a8c1964350027a8081ee99a89de7ca7a5d16360936eab5210c1672b53fd52cea6fc6286a7cb75105d56a744cf903902004ff413146132768b5f004c7264b1d69cf6fe3d5fe4ce9e7c18931bec44f714a7028bbbdaafe3b74b72ab82cac084c8a7020a947a540eca3f4e2de3d6640b249aeafc178a3e7726bf13b4934d26e08d12fe017f2f75ab010da1fba6abd2266297585d342d9d99da7eb8465535072647e237e2cb69532352cfa6b1ac442d57e408f14c38f5a94cdc46b5efc88785348846e754652f13b214a17a41a7c5fca0e61dcbc24101fea1b393cfe055e74215b0f043a1620dbfeeaf88d7d0a5f6b797e9bffaac949b574bcec9552bfbcc9b1a377299
