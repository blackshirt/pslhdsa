module pslhdsa
