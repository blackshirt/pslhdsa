// Copyright © 2024 blackshirt.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
//
// The SLH-DSA Hypertree test
module pslhdsa

import encoding.hex

struct HypertreeTest {
	m           string
	skseed      string
	pkseed      string
	pkroot      string
	idxtreehigh u32
	idxtreemid  u32
	idxtreelow  u32
	idxleaf     u32
	expect_sig  string
}

fn test_hypertree_sig() ! {
	tests := [
		HypertreeTest{'9f86d081884c7d659a2feaa0c55ad015a3bf4f1b2b0b822cd15d6c15b0f00a08', '00000000000000000000000000000000', 'ffffffffffffffffffffffffffffffff', '1feacb19619835f0637c3252d68ef7cd', 0, 0, 0, 0, '1d8cff94837952216aca752fad2bae148bd351bf7f72e44ebf88a54ba30621392af92b1d6ac4d8a7425c2685ea6c47c1eb7077ef9817fff78dded68815f36dfb9fb132d18bd833ccfd093d6bc79c9c9a7b0b1af2b88be036734af0b2d4a64ac216e64cb68f0fa075e12b08f1370d5b2a5fd923e2ac43d78eeb82430cea93ae398802b955817e67dea5119b9e27b7eb30c863a644371fa98c275220b16958a671cd362216622b840c2821fe0000f99670d6579c2a604d85d5a4db21bb10784c6359dbc5bc3ef3511e90b46c5bec9c8045e52d6dd25c7b04f0231288db99ce04adacaa3cb1a61523d3ac147a6563169f822409ff673401710ee8250c073a0656e0a35ec35c6dd953e52141fc704dee97d3bd04e9855d04bc37d792bb8b1e60093c802c2a08722d9f9f90e5eda00448c7fa82141adba465b955fd971183dd008d26ec4efb8235ddff418832e073effcb50502d7862df634c05aa74ca40e854e4bb5060de58d0e479b941dba4452eba052f88846494e2a6a1cc1046ae2e26e9bc36a438fee4f15a285d09bb7f17080a9e62ab6dc4d6120f014bda703779f957de6f46675c1f11920cfbd0a9b2b817d84181a78f59d3d78d6b78598c11667edc5e667762d092a1a6ebd24b1b34fd37c7487fe879e2e0a1e66ee99d9e3644432824649a0cc4cf668b30232dc02167e6d74e0cb5800178438bfdde4238a05a44f9031551efac16d2824eca3294ad3e5468612993d58cad4a272b401de6764dbd06f09bb80b62585d5e1944fba4919bf697a0f92ee08e6ccff9f9ccfb7367d0f12208c3ce1c9b0ecffaf10feeb754629eddb6a9bc468a4f1b435830f6cf3b3a399b710fd63830cce0d7fc5ac8f47417b94abed1414311829883510435fbd826d958d99f9dc9e09cce9a2971aa575414cd4835a4968d2eeea8afeebf1d249b50545760aa560e2735e6a36b263cd2986fa9f17483b4c2f68fd45acb4281ad399fabc7cc9e2e66dfcaf457ff4ca89aff7a868e8412d685cfb99aa92ba14db2b55ac0fc837166b2e6c62ad1ad8f28d3be91c64efbd23353e1ddf5d904d3f63f9d653573fb23aa125698b44ba6f10132674539e4ea15ec380f2ce749523a0aace9c7d53811677407237e2e18b4609b7da6d7eeb163b60a4d14bda1d7b38f015ef29aeb8d33f8c0ff4e2399a1073ad97941abea1145edd1537c3fd4d7c1580b72e3ec71fbf44c7d3cef3c6efc5e7399a05381e418664790ec86a65d5a1753896d396f9997630e8503ab9896ec9cd31861b47bd01b59b24e07a56862dfc450601112c0d61cb20af2c788bd8a7097193038390f646aae7cff3da22df3fcf9bdc2d3c3d67ed384683016dace6b7ef31b356138aa8dd70acc22b32cae13324a45619c2119f19db98721931da9767ab3c0ebbe8d9fce06f109097c7e72e51b03b62a408c6d364084aec922da0edf75040cf00a0615f10fe171d05d90cfc3988a2ec28d0de97ae0f9d0312652c1b2a1b418024654f693441f6bfacbf41aeae3bb9db6d982e04354c4d135e535520614aa272794cd7fbc345cce13507a100b1edd856a2b7cf83b7678801b0b6e6dcb21cac2b279b5025adb99c5b0fd0bd01fc75aefc75a5404512c5bc4daf29f552d7a28c973c51f0a71e515d3bb836c534ec51994258bab41508084a4107265adc67136522875bccec5c77e42252d5f03411d334a4e0c9ebdc373fc0530ab4f361b6d1fa6da05de631dc093323a1d7b472747e2e15c3096d34c7e62f4a5508df334906971ab096d3f069f4306c09fa811b7714419020b43f5866aa3ae0d811b7e761150c95a30c42e5b59fc606b24ca7a7bf542367e92eb1c12c7ee062085bd2ba53fc3701f9328916708aad4665f4df553d6123676abe98ddac34c1565a75ebb1e28550640666472137b48515c841b843b078d2e8caf411eec2da78de0be1553e1aa31ecd21fcbe09a873558fdae0c1510a935759390c5b45110bae9403bfde5d52ee30702db90bb2d9f0aeea012d8d9f1ad700eec6021a0c725b9002b3b852b70af45069f5520ca8b139ff916b49b3eec84a8c8e9ce33192270ab026b03bb9fbd1ab800f28ed75e9dfb78d3fe2f482a62339f34bf23045991d0034f6e8d5fb214f7dd75dadc7c640e2a4c525b25918b82bbeb1deebbf3eb2ed7a522a46fd1dd12ca5d10b64e468d2d2d70e78e8342e4fe7e48ad298bbb83fa1afa1c2d44a04b7b08688dce39c9b1be4ea44ff2b20709f03b8500aa3ce1950e9d4aac50ba0992f08d3e389a31ab59e375278d4ba3045672d2c4ce85c007c5ad5a075b5ccf1c79d12e0778c52cb4b7753ad740e409705decb6bf019836fecb5b95295180512cb4b2061f13caf32d57d4b88a4e1bfa69564a4d478c8cf92a4861ab2884344ec09748813e90b792117a1fb359e87ccd5be8e5e4aab2fd36aa19cd26cc46dba1a1e0a1ece8c82c7dc61f9569eda59fa06f999b1ca796934f493825feecf54473f3cad00a202b0fa7f29acab619ebb2fba33a4a06a9d28e27aab775a85b0a4639a5fc073e898501c0747cacaf65fbe4db06e95c0d6fc6ce33f9bc118de4176185a517ef19eb6969e5a08bf4bcb23d567e4f432894913e1823c01be6c5dfe53539a8e142d4566baa3cb7dccc501468cc3986156eb4d05afd5571452ac93fb80f70ba8bfec971fe9cadc953d2b80aac425e09e3517a624f07c8149c1961c0fc3b7f344a4e034b0af62d8470412d891a01a0447e37224277fc762fc7ef324bd1a06a3bee60be7f39e39eecc74b2963e33c29d22cde29ca5aaf68f58a2b29c7c10cd8b8a37a6cfbd3583800a2832b520063498c98d59587bf95a4167505b2cb67f66030e797d48765525af122b23f29ec41df83daece4ba0b037a562e3da5e2263624a3612b676e3d17bf119a615daf32063fd14615dba5305b2cb294f25667fb1bafb43dfb6c1268083fc0a07e8eeebf97e82665429034053e560cca5da65e64390e26ca97e26ac08e97b15017d47c6fb8140e3b0dd3f9de838870d767c47e0dfbb46efa9c641ea1923d4099aa5c5444b68b95cdc142748995c1bd1e80b5e7654073ad35d3c3b6513af5d157bdff28133c658b9291ba828c9f5357ece2533bf5a7f46c95109a54b6bc3c7e6ae78ca5f8765788d8073ef4c71bc73d9e154448090f5e0fc28ee23265237310eb92aed2cd0ea66a66fde66dfff49797fbceda3b4dd30baa4d65367163970dce6408d20bf8acd99949081381badd57acc12db8c33eb19cd61f03c00e8cc08cac5414a602959d0765705bc669bb648fba83d00e878770dcd07e787446355fe9c32cb81104922c86f85d108812e95122ac73dac1ef3de295564e35751d920f421930b8b29f525b06593a4cc7fa180e186ab69f1248293869af9afe139f261f3fe54d150537388b54befebc16c06f8baf63c8fad6cb286f1ce5887a697dc428d9826d445306272f649ce892fd4af08b3215c615e7b0c4e9af95a0b5de34849c6eaf3424829ab5db56f7ffe46e34d25557bd3100e61e1b1729709b26d6a8176e82491b8fa809be9c9dd4719ba4edb1c3e7526e4789764119315dd1bd9f9e5845fff0d8c55ba250f7b8758c1cba9089e8f9ab51f39b9b415e52bddef804bd82576d0bd49e2d4b988fc30c1e3490fbfd246a547ba8689b4e277aba3ef15b926b0a68975958545f750fd71b4b3e8042cc212e61e97939f82c45026e0fcf805ab3df557297c1c6d2aaf0900f56e2318060cbc2365cd00e9857b1d5a4da91b3aed818f43ee08723a2ac0876a60e9fea1cc166461c74b8a94353b51cabe9767e3075aee8f3cb85a9a43e24d0d833a77d4cee0e3e3424b4d199b2ac00ddde6ab24752c1302c3be546486b30e5205b5cc353b8cda5e0476ac10b066c20429ebe0f6c4bfb9195d38b08fb9aa21b5cda8f01a763e2dd1e60c9a724a9fb05b6ffadffa92c7d7e33ff8bf8a8fcfce1e33114dc4de526ea47cac6f7e507b8e519508089f5547879cb94c8c8c1c26e05799072e36d412f05e2168d17d895a516c4569bd6af198ac46b711ff1d5c5f53c132e4fd5afa6292074f38a633e277a2237b8d9c2bd97272742a49a210b634e0998ee4d89907019732d598a8563d63448544e467727f17ab03130a77fdd07f38b386933bf77fd35962340faf8ec9b81c33e3d79963fe5881844ac4f85621c6eace496dcc59b05a7b824d7209866775f131de79092314c16c65f34c02e97666629b51af98f7d4c2f9bc7558d8917bac529df1d2154710919a873d796991a7586341db7a7722165937659cff82aed7dd4b6252d775ecd37eb92df89a5ea087cf73f2b53bef28e17652d25f418cf35cefae37b9171340af33b38ca5b42ac5a2916f7d92f2d6d361e0a136486355b2c8572a4a6668e2ed364fc1ac7ee23d5612c5ac25ea5b6e07792d79845b6bd417631c6d4fc4e3dc82b57d01748c5be27f891122be68c6a03717f3693db68ff465758e77a97d473b21bea4c8f026f48710d80565ef36803ebc908c08b7ac252a9a19879b16a0f85511bea1a5bd7cfd983a519495cf16f6ee00fae5cf4cb324c8bd431458eb2cfa86cd41d8cd064770dfc56f4ac5accfa4c5a4ecdc029997f6dbfe00a9edc6d1740a6acea7434decfd1f84381d529e98e77d8cca6748f53162232329d66238c08bb66a9717244f731614b0e4fc74aa64fc350b56bf9935c692d4278c0c27ab9a08f2328ed4536716fddfc653c25a0e72a7ae00ad11251c7ea7e315eb752ce9d32539cc18757ce74afdf674a86315770d52b6f57b5755cbfddc7e3d0fda5f6eecffc618b2788a2f1a4950b0211d44226f84e8d224594f7645d50cd5a06296d50f0cece231036aa4b60bc2ef8e98b44869a3d4b7f8e030163ddf96962eaa520e522693b8b165fd933b7170537651bf08c2a35e26fbf703e536e45649a6a75a0d2cea057f7511924458d70f554283b1f319377f807d0db7dc5fe400f8d9a3938c79ce104e65764e97810ec8f4e181f069df374d7bbb38134f37bc614c81756179667be33b0ee77427be64156282e8cccd8f719bcaa897efbff7eb3395531db81261f892c90fdf6aedb779f2b2315523b4ea79c0a7068ce2fc955d438f57fdf01f7decbfa2d41d1357ccc0bcb699b452a9042eadeb7e3a9cdcdb4ebad3c3c4ed124e973229f73bf5480176403095390bfc6c845a6c3d7b8321b0cb9d6256baffe3e3c1a396a44f7a4f81d3ac6b2a454ec7f349689668fa4facc144356a5e545ce6614081c3f4f2c94767a2b2813aa59d703ce6c71d042056ca14d976814864236704cd1ef4d781179ae93ddd4c798a908fe56c861997f516a21bae89c2e6a5e96c767ead3bb1fb4872b4ee6a94e1b26365d9cd8c78fee91a939ee5146f1b5a9be5f21a2e448e82e695175d206df398f02c0c9577de0e29c150d08f120380374abee8025ca9155508b247d1f37f422c7bba01ca20693867b5a040c37963d9e8e787d537fdce8f61d523a58cd6486f2ef9f2ad2b33b759922031cfaba060a43772f054350a5cea5b63d168b92cc5dbc94f527b5fdf694cf1dd32d10ccf9797a8f89f9c30f646050dac61578148a18231da760ec84df9b340e65bd8d36ad0fd583fb858d2ebf82c5ca11ad372ba6b5d68c93803dfcd035d561ad0dc28365b4dac67e4d958cb002f98d889ac0236389bd88c31fe3065bf293963b94c7bf327ca6bf2876a673a169f3c47fff83dea1b269dc55fd6296a98b990f3fa73c3f34d3489ae54fc430549a8b4dff3c166d23ed9c1c94d589898621e2f0d8f86bb00e6b1eb212b05304ac5ac5a312fbeff3e40a1bbc63387bb8f4bc12e8b7401fec165752b4f6b9abadba10cfc6c3e58eb4bccb224f7f047d304b20541ada809674738b88b91dcb66f671fa053e3b7a52e3bd3f2f2aa5b182984fdb92dd3e0963d267ede82a6359aae3ed1cbaf8eeff3ac354874d4bca2d5c5b3291564f05468bb7ee3cf0978a3800c48c7edf57b103def63a9238abc7ba23b26c78505601e493e9ab0204cb0b2f6b7d596c800cc396b5700fa5f7e45f8da3afbea7d625e6455619ebe8007eeccc9bf37d90faf40475eb6924a587cc1697f46808393058f4dc8fa8bfb2e2e941883256f58db7ff6ef97f96b70c8df103e9603fe813629dc389a6ad615600e7eac767ff2b3876edac5da2df8a3cb39323c1e606dcf74f7bae19d47b33e32fc2981c08fa717965e09add84065e2e37ba47cd727da01ad279af2747284bbd8a47a5c30713b8b3f8b6e502ae0c3afe0474b009bc8a18ec177d0a952605437469cc0003d6ee61379446fd9b391333506d09534802866d7739bc7c5bf098acc6ab41a3a5bef5c1357b5993d06d7518086a92b80b366e843405d4f2adddd26ad6346e11a0fdb0a2a95526e6e8c588dcfd2fcb3aeb3d7c58e8a1ec02ee3182621759bb2df0126914283cb613222677c3ad9c7e4c8e9fa342b1e2c5f5c79ece196c5691b83c85b24a8cfe09ee8a655a6449fd7abb8a8ebe8bf07b6375bdc66e7845d483ae6fbe2982187841aeeca74c8ac1ebc4343a5e8d7d446cbbb35fc95818c28a9edb8b56cfc7723d107d63209d89d7922211fc405be3aee70aabe4a62c4986f3e41c88c6bd3a8196fd5f54aef5c76e99b0ed2a03ae235575c563ea20058dbb15fe9c92261276dd50cd5053140a3370620c99afee2c100ea91f23d0e3c9f3b5deba7cce915e24e8ca7fa751778d4f23e94cc3a96a35bed6ef2b11912ed4480c8645991a56c9933f87007df6f82432e473a25237aec574dd3b3f2d31df2d7df01d27c779d212ce7840830baef981645f17e5fcd545b8705d9721e31e9f387016e3f3536aab1028631347d4442eb050664d489643f066b9fd83a224aa9c51ecd8403151580afa0b0b2ab80ead77620420bfda1423f4c8562a657fd7b82b55804fd5f87926681ca1bd910ce528cfa487de482e44e9fe76b2da934393a3f06e3bb50df9d9561436ffc77cfbe11fc053feab934bcc6422834c55edbfb6afc39431f1ef4ed79a259412e19b3899572991693a0dd70bebba3ef25fd631f076284febef7c6dbe1da203f2bcc55c6d15e92d4b0d167f4b4aa7bb0e4e54d7f6cfd18f74e3853656886e4daf5af6b11f98030595d150283d1aad0d32404d20586766d63becd8d5dd933658e21be0c24d09d0c7d94bf9c3371906be1588bb23cd212e6f3c06a6fe636073234efa28701177d7bb012e80cdcd55b28fb23e1c0a6f7ff1635adb6fbe32e36a1ebcf8af13554a3e70de6033fa4cba4bafb9307999207dddaf8f2fb88fb4c0d7cf07cbe51f5b8189d8c2208faa2e27605f060350bc2bea351b9b7bd81eaca1655ffb7f9d37cb68d5f31bfb39fc16891cd85b3c9fd9a90dd1a0facf2a677578dda5c9357c56960c078a2b5f02686825c0726ee1b7bbc1534cd7d8dcbfcb2283d4d6c7218388def27db4f4182bb149cede23d832596a0697ad779a6aabffd091ffbfd83b2d1242da1f844522cdfd7e9bd404e5f9aaaaa9113788bbbcc03a58343dbd9538d05cf4006b9a7ec2a46b2f3f81cc7eea833f275a83e68253243b818b1d34ba286726ab794d5983dc5e48aeeefe85e68f869f3db53d699f8bfbb68dadf032567adc68a9979dc7676fa2c347f3f766e2f3189062d79abcb51565852bb25e51854f73dc6067e9b6d31e66b262c002206301730a4fd144a127d5ed03a7ff5a756bb7458e0bb42387012bb550fd88c837946021f84615877098ac37afbdcbfcd938f8863a7cd4006c69e6c6aaf7b7bba2045ef98f0ef9669b657c128e5268f63ffb5d55b76dd0032abd5e2569965d63f30a0c91ce5deeb774a2bafb800528778eade032a0ab1a389b47a37d767ac5098a150e4e664b72731a52c89605a8f4a74b40ca7fed56e8a9486b3de8aec798c593bc3ecc1595e6cf68a6723e9c9c48735d6d78346a5c1899b37b8833830767a8a8fcdae8d95873a9810c37bdbcfcf93ace21193fcdfde3df6eb6df4aec5baf4b7df88d1e3f9d31be267d6d5a9e30fccd68ed855d6b6157f58e3c478049c5dbac3415832854ef33e3fa9fba5e51fc5d2afbd0e3e1394e189ac10d40c8ac23e03d4d83355cddb4e35ee3ba1a54396b481db5c5074265699fc5e0103b9e389af0eb909f75e2a30ff1afaf9dea2015f3da2f157a179a017ac23dcb88f04c0470fcad70dfc3ac2855ee1fbfac493afce5de496afa111c458fb887f9c1afb023f18c152152b464f9e29970c2604e9d9e4157caaeb0814f6694857d9ba596016c3fd02d7306f707a9fc3b4fac6bfb7bdf1ae287565c806404fd76af62701ac48095459ca28f9c9df5bd9ff4ef6ca60fba398a9b3411149b852c2470f3ea20aec51db5ab56a51d8743b0f8a17d41ff0769264746b015a17b3e513c504a02b726841b8baaff993fb455575a79914fe12ec085827f5eb0ca2f459356e58649d010f47e094e191c9d6212a38b51e99d926a30d8242bb20ddad0510e799d87793bbb2b564047688b85d8fb0491e447874a06d12eb415494c575c7583aa0849a870c386222e628bb1b2e3f99c098abef6d009275ead19608e237b71fc814db60ca159503c8a20e3098151552bea31b36969d3c31b2fd6aa4a17515433a7ea2b5b83ed39fe7fc2c6aed661eef0c91bbdb388b12c9b2a24af59179bac959d8532b350020fef8c6b80e584db041818c12f8a90b9498037a3913c334a4877f731ac2e24ca5b39c660293824437cd28093cb1c6243b5765c679e616b0163ea444e7578821501ff69593a2f59d1ec443d82ecf1697aaa6353cf223feaf100819e1899ea3b0baa29df19d36e452a4e98a7f78fb4eeab6c52998c3da4af83056972fd603a1aad0a8f81b4253e1f9e2b7e8ac835307f3bc1d8fe5543af1caee18437461ae1b51726bc41f516fb60b9ebe789bb9630cd2b36ffa4f51669053d3868f5af800b82841e1ef586bd9981de67705fed342193c9461a50bc339e67675efb4d4903f4ab54fff02c385792b287954131ed82f6ee7322c4b1f9a58894226d3802975a1aaade1119815ca59818e45c7ca412b7a35ef7b4d520c389793e2d2ebe6435ee6aad09bbbf6bab4a1c0a8cc135ed55221635f2178c5ac78d81f63e385c62ddfed731f65a3c7ecf4704fd3680401bc1fc3c135b5ebcca231200589133ed38a1343427d757892826973f8977f6306f1307bad215871974cff9209eda611680ca2d3c8ab29ce41f8c9b0a659b26d507cc25755543c1388a2a525a556cfc87db08294af5d8168158bbe5454ae895cc3ad59323fa0361750a1bb9c05b1d37fe41fb91ec2dc57347dc25b81fe962ceab821ecd122320eb3de50d9f10f20de99d5335d702eff7bb974c04c2e9026cfa0794f9f58ed9ec513af9a1d5de01f09a02e3b9250754691c6ceac0e0418e8f82289db8e8778a5671b16f11d50027441cd169afbc9d13997a61cbadf542fc8b53cfda90f8de076f6425e62ea8c899b3cc76969e19dd494f16a3c817f7cd33f332d0965857943a36478fef61615f128181bc87774fc8eddb63befe56964714fa5df888992f5eddb1afdf65a0f1b9e8cc347dec3aaf611f2d634f0415bc2a739840f04df89dc3defc8d39fba9168ef021bfa31ba0759f6a9521936c29976f3e7580ce3194593630b023ac1ec6417e8f2b3300b5cf03450659056c519610d881f81ccd487f24475fe56f1a3923332ec4d16fd648821dc19164af8515a53941f943b77891b0bd8c695a68941b3b34cc6bd6e636c2350070246234560f763b5cc769be3f59635ebd487df9e9ac81a6ea8c07ce865287bf2b9c1b17e639d1af681b95b6d06c0c37ec237a40ed0d0c14725f04760d6342ef9e68f99324481aa17368a5260f0e195af1007b6cf263283e0731eed0951b79120f8ab57b0d389c53dc11dbb40109f34dfcbd6c5fd7c7dcbd7427a190911a3937350e23050856c6de0b8f74f8e5157170fd1c2f8aa91008d1c4d7854c0a3fa79e4377618ed4dd25c17b83d25a2ed89310076b51d3640d621deffdbb02c7baa8856081b09bc3d001db2e14be2d73d397cbb0b9dfda73ff4bc9618e13b89f4a05170980be416f1eaa7ab054f22d8c4db28d801058d940eae86a27c4c876b23b3e101f1a9d5762873ba4c2eca0c30fbcf855a8aa895bd5f0dbe8b1452e157a3d6e68353e41cfe39fc77a156048034c1e68ddf950da3fe28fa613c82c6dbad6d72edcafb3b1376eadb2ba49c9fc34120af036a5cac38a8375fe5c6ed1630fdc154ccd12ca85b49ad61dbf96607373bfacd2b17de3225e6e6a92a505a9078a0fecfa06864b2e8fdb4a7a407df49ac743350e6a0382c9c4ae74ba062fe76b3e8fd8fafe9aa9df1a3b3e288232f29634cd222c06e809fc09c2f0a47d6b78b93e91ef24d8ef0218141447c3b45076b09b69d9fd45bcd8761213294c5ee1a839f834c7456e9db336a8326c82b158c0b9b60708c340bb5751425dbe09f3eb69882e44b357f1a6a527e28b7fa2bda0021d8b0e4c0d850e1087935b4a821420b8f4b11ad19d9df18aabbcb714c4eeada962d748c381cb4e94d7e4e93d703565fdfb5ebd4344a278a045bc7f9c766c9aca3dc4b1ab00ac01833195ea76d76683e72328a77fb37254c9c3b22615f898f61dc7b7002b3471464795ceac1c55aed8540777fd2ad4c65c61f3febee1523afc198970efbdd16eb5ef132a1cf3bc3502abfc2778281b03e62c4283fb84ed50dc578480c9b496f7c3f1ca8300b49138e89e18b6981ad04906269dc54c5b48b97b710de9db2acac39b97eb991e10ff2e517ed8a4432a48447ebb50892d332bd6ce5e4b38692ccaeebd7ab72070e56da4d946b610e74f0a4e62d02002651bc3fb95bafaf2802d8267a228aa680afb52825a9aa3f0789495be44e5dc4550bcc0510e0ddf03e120cea404ce747be41cf20536d52b4da9faf60b9cdd606a898dd0cc4e87f30b47723435fa400b80cb13a1a29501d2da6040a4e551d6045a5d110a05431d2cff6b96a0b488ea7b53031858029ac896d3f8a44b8fd5c5b43f34e89c093731302e394edb1430a232174b7b52818d55bdd9d40bf11e1bd7cc7b3a133f50c9e2693190a4c812cabb016c827d92f1cd6facddfea7f1134ee86e0e0031d0ebb777fcf3f35c3ea4ec0e94278e499a0f76171ab9ef87b4249068429bdfcae641fccea914874f3c1c865ea7521896f302f3e7462563e406539e8752db86dd90dfc6f7e1c3cce58a44c29e154e69bfdb8b3cec9b84ff83196f550bec78488f63862541a767a62fe4c883feb402b0499eed7aab03e47d915dcedc32f2240dbf6f215b59e6ba56737556f9a8125fe0e3052265c0a3861e72af149cff712b391e0fbacf5e943481e4b429b236c919a06bb1ca986965917ce419889d083280aa13bfd3eca4a8bf363e31bbf0c9e9951da2006b62aad85e0e67606a181eb3319571ad7e024f210573ab2715063cfab51739e74acc7fbdbabe4877d5bb697678527251fd2c445b44d2a079a1f97a274ebd94754a8ce12898ac5cef9dfdedb933f5da4bcba79ff834123b6ce6af8c15f0b6f798a7a6e331d4f6133a2e4fe6ff7cf3c8b8819f707ad1ed95deb1c96e4832c1a4d068aa0e0ecbacc37a01d6d823fc39750e765618b90212ff248dfe0adb99fc7a616bc299695a2c91883357e6afe261455cdd31c41924d34c0f126c6e41197930ef8e91f1b91bb440b829b56c9d6a2d47a877503d3dd1a80df9c52e2ea119ee2b18ca88a8060562f5e28fa6b934f472ed6757e084d7dc9222407c62d556bfc43dde89918929e0df8a4bbe753b7b1268be42d4567851f7278decc426f96c688be4bef6a8aa90271bf39b75ab734459603e2050855082dbab315aae0b13ce61aac570a79c127413ccdeff786b5ceecd84ab2932e57ffa75d8e2e8443fb0b3fecdef38bf71f2f605eac1fe6889c82c54b27ab9721c7c200f61f6f8b627d7304312bd4424a5f25288e0af17f3fe3651855631c2a4fd9d82f4cd4ec0c95f92b2ac9909ca3f20668c2881046508a9cf531bebac970ad4663256433199a5c300cac62c4f3af8652aa10a8876f485ccc41171f445c9e3d57eae6aab707cd94f3df628a0890f4683398a37079dbe013a07952407331bba57855057acdd9f7b283cc71ee45c6b857f519b34cc028e5622cacfd0bdaad8a355590a30efd27ef803ac2e6f3ed756be81b207c1aa9e706d4ddd142c0166975397b74197ab4ac38a1b47044cd30adea6b1f7353c3f5d2fa28764381c0b576b8aec3a49b1727dcf387b68bfcaf8ad02eaf5edea2bcee274cb1d2948518c687570e9e6b7ddf6bcc3266497829c4b5a804bbcddc3027f90a3bdde18bee3c6587f047e0ac470b614205d11d127558f369284cc24764ca22bc1d79f14f7caea3d846d4cb51b0477cd8f6873b9a3c9c186ea0d6c22e2f9f8ee8da9337161df74659dea26177b27857273b7a792b88021f68621c4d293be11e4b9ed88e69d23e60432cfa2bb7ee522bf2ec4162f68f1ebe6b07b0076acafdf9a4a1c26cf725809dcb4451eb5d404c7f1b0375340930690c10435208f446d7298731ba7359cea724d1075da3efdc52d5404ca1bd3135e59e0218dfe9d6d0287b318ba04d3671f38be778402cc5f17d0eef3386a52eb3412db3c4d2e385dbeb8184098d7e23357b7ee82ed59098ee2ec4f0316e0c7112e8cd2de8e6f829cbe2e6060b2cc776eb6a144a20f3dff66a94090823abbe80080347f2de46b0b78a98a6d5c4c81eb362f608684c92bf34a61ac39d30a838bb7423b40f6838a2ec18183c098663282c4a9c575b70690e252d07ab58a6032cf41d3b41596a31b4caab82647d53cbad06a913d05b7d3ffb13106033f87c31ee059e851133868c88990d96293d654a457c48577b542460f035b4bce994b822bf5795c1b28a8f57cac4a1b9b5555374b569a2a9005657ea1ee492c2bd0d196632b3fbab1526651cd1f071fc63a918b6e3bd09101b28205f53627030125401801b75124ec04fd90e0cafb58e3c6745bf390de6fee88f66a6b79f0cb7b8806b545622b4572151ba4c204f467a5a8399af2a401554fca48c6c834dfa3ba026cbfd00918693d6c17fbdb07d3982bd4fd6a17de1f94f211b9b761a05663a4a4445c96c252903133ad73f79037e1c1f3f11f88cb25d715957b032c63a10ba4233f92e3bde0f6139948cebc3b45be94ae4b547a30aa42c98ca84d6b235a2b2446e97748a3db7a6ea837bd602806d9f2825d42cb7304e46b8defdad32c3a0183269d6419b4858fc98d2a76270b63ec2af7801f124b8f93371af1de2afcd0515a576fe3a38039b4d096d82a17df44ec945015e972729dadff4c4aee4c01c0e77a51f80e9acfcee9412bb9824776e781d3792fb9881af2f8177463790e5cfe57f4ec000ce0b91fd7a174826235036c369dc6cb4edf77ba1298e68abd5e2d1a1bdf42f3cb52674b7ea76a8365f5c6ce6cf4ae64b909a97c1641e2e4473fe00b8a49ae7cf382450cfe646448587001b0049fbcc09a24d47bd9678301d00b4cb9e3958a81c40f4505b0aeb8e768087a3e79b43f2f2faa5b6449694f8dd03ecf8e06b1933d8cd042fa8d19c7b83b520651657c7e8697771f3a6689463aca1c951f902f7a799988112fb959f4e453ec35b4c1f8714fc6611944c09ce362a0a12c50d19301df8cdbf8b8a247179829e80efb266f533d29f1e1c40643f5323debdd9091c87dbb17d7c6e9a13ee78026283168ddbfe399a842d4bf8c219bbd94995f46119a98985be217db6db6e11b6492490a8d02e3178f1526beb5c6db79680881a6f0c1e37f14cd70c7ac26650cb680d4800b18987c06f8276f362390de833c301637729fb66db3dc15ad7abebfc2669fd29264ed14366a5e60e3c34b706af36f485d3efda14c20cc90388d99f1a8b3445b415c5379e0c4fa67012e28eab69e87969fe75e27e71afd6a91f4d3da7e2d77f49df66220ddf548e4bdd16c3e77f562a8dab02494b9faf8ec2176a46542c9e6feb86a1f4ca9e3513957607eaa036fc811a5936f4a8ba4098b1d134239425d1eb958f90488403d6145596ed8b664f2bb3a5073e15e32dcda8b10188b4ede8c1cdc83d61065f7942abb157c5f8c0b1066b64a1f094f580aebbb3ac1428549957dd0c09697dc511f17fef38d7565c7f1f1aba8a730f68b39c18a30cbb9608a451bbb7c9cbae7a64338d2e6c841f78fc43f11d62a2e8a5d61ed11ec84355cb52a64a2fcb74537fb50b0c15e86a534c78aa5bf22e8e7ee88bb1376d9e5da08511c01b02bf7e13a8232ce1e924bed86a209838f6e406ffd76649ab16f8eb39f406bf8bb57ca6e8eda4a9e8c8a3cdeaf159abfd3b3f93573f32e8fa05e0d971627796e0a2e4a4c9d406fa91f6250a702a03f6c243e8b1c15f0a6f093b41606382e5d951270652fd051610f787e4bbf4ce584a7069373e33cb25a86cc4ddf7c267a1fc73d98737ccb57251c44b2713350785c0fe62413fd69b724cd38db1bb422c338079a38ebaa4dcab2588d96480360340d290b94c23e68ec3130a205c183e3c04489091fcdea390e8b4dc1491286815894d36da7e1b50ea1ee89fbf6ff348c9febb799ecb366c19b88a0c9fd437a8eab1ed9d24e616de7c9df870f074803ee0ac1b8b354afd25703a28cfb17d7c7fc3e214422c45036cd58d83353ff24bdfd76f6794ca35a5fa61ba8fdd6566819f736b3a21bc0f34c877261257dafafd8fca1410fd52c43b77c7edcf333db3bc88fc4ff601f87304a8fb03460a24b4bdafb271bda9987786406fbd7da368471d095e259a800c64cd53a57d506a8ea7862b106f67a747f8496a7ae37870cb314defb685e55ccfeff741bde2b335821c878b8ba16183bafbbb8468338f176d2c953373f4c6715466011d4b7c3efc4068016fd10178e5f9e03cadc48dbff9194d204c6d9ffc7b193f663c346c70ae452099d40a73d77247c6dc9eb17a79d3a306ef142df8926635f78e9a66db9ed565a09dfb845aec1646e500493b11574fe57fabe1c68869bda9c7943a685253a5a5219fb7200d2c7ef25df2fbd053cb55d4c19e30be545e4199be94512c17cad17b5bdae76b5ffeb9b7bb28bb880704a096c51095bab729f9b97b56818440f29faaad31d6480617a8651ba245e78a4178cce67f0d8eac91dd80dcd3c78c5b1a05800bec7c540174fd7ef20d5e63bf0bf3d7f15eebdc831437cfcb016e2394d2a8ea7cd5c12ccbcd83f862ff077ad2008a0c96ef60a05c79be70754067ba3336b7b96f866e0f6ff84145a716d2737792a239bbc513aa26488eef8717fef5febf28546d7671ba6bf3b6e199cb25e85c2c18249531a206ed5a52424c2907a2bb4acc05a3a62373bad6ff0e811d658772f3ddea12ba2273c49de28f0d8ec08f8578dcfd5cbd8ce09ce4531623d6e5106be94e495b86dd557a767368b1ef7193b52894cb3de048dbef0b2d4c5ac9a0aaa9f5ef3fcc620e1dce89871fcebff669062889cc10f1a25d34c1b726b0e057cc61a18f6e80dc3da2f39a2948b2c1000d0097a6c477983ce5ef0d289adbf2c3b4e2338be49b61a9b895c2a9729561e4fc242f07420a91fff8c8dcb6219a07813f183442c3b4d3b35c833d7784c57dcf77d77c7d03a0f06472fb307b72ad6c50db78d711c980027ee113c5dfa73ca84c5f05a510a30f82f7297843368dcb1aaf237f779d7902a2b2caec9d25fdb5ddf24e82b05a54a2188aeaba7ebc8d14af0cb82531352a223c13ce6ea726983a2c81a207a2efa7d29df8faf6497e731f99271a85012ae4b95d975e6245db4677e37378797253ae6b054b879f6bc008e8010d2728bf7441a06aea785e59b5a5f5da424bba97ba83811d6b4d2b45bc8be79bea0f20d76bd9648fd0540aeaf71b1fd2c16854bea8d54a2eb388be117851cece668a44b30a467e47a21c2b2be46c36e4cae783d2e24a781735bd12a9e21d8fc5266e0b872dfcee6995ff42c50f91ff5ff4a59476579a0603ff59ba6af2fbf67e950e88a7307bc3fd241152515cf08d8e3b51e0be0a229550aeca37a50de1e8ca4ee2420f3ced93d842ddcea5dd2e8167cc4c4332cf1a59dcd95cad9f4c83ef6032eb4b6ce9046020155bb6bad5ce3781623e2256d36b385625e9b52cf2e862013e3c71f848819f72c7aaf40a6215beee8ea628e30adb490c65b225097a3438605706216c9bfdeb11046ef7b09f3766dd2793bae2f10127c04f7a6120a45a1c5c855ef992f7a96977df00f318c2b3c4444119881108614503e749da3ad19a0a5d00ac45d406a8e882af7d3b6d584c61bb9e3c81c8f4daa565a7d88475cd98be60d07f3247e2aaf37c91fc9ba3a2e84c2eb8df2a46ac95dd04dd459c600a3f7748fe5a140592c184a78a6e79a8a020c9f6273f877633ddde6f735192d46447b090c16ad7a40fe0c5b9b4d95d7ca90d6815aee2207334f60e2ac1b5aa8db12ae609657d4a679d7e4529116806be25ef5a3b42786fad0befae4546ad928788ae55c1226040584f2ebceeac703f1ce62e57d9905f98eb06b9ffd77a2ae4c638321166a4a9275e443f76f7a5d2e08f3b46c18c62516fa84bb1c82e1c41fe74e236b7d66a4a8cbe72f3f510a4e02b9100834a5ee5765e272d8c26cd6bcbd0a8aa3d33802b86cdfc9768ff5bdd8661265f3c3fb8525302837e6f5294bda3ae3346c5ee57a83794b067bc7d844d5c09dadf7429f09e289fd1f3b3542c457df7d03c197886c35bb29fb8a0b9aa2cc68e4ed273be91224ea8fb97c0f4f50f2e867c562473e7a343de6d3796ce91ab96b5687a2fe1ad1e7ab68a0eec3adc82e744f4ed6a935c6378a696eaa8e735217cd509daec8968dec573d806880c0b6548aef839fe28f9b329d2d97f92ec9553ec1c9b958ec744973f314252a00386a7a882390a027b2d99ab295996f3d2700459b9f8d4bd9c864ff7d471cef2822a486b35b58beab281cbe29684f7efa94629d8e4fd706b47711014db840a72313ac191a827cb00ed0f73383a4952e72d1a0fce1fb319b2f68eb6e1a550d83622caa855e830d0e19d0cf778c8b246ead0fca1f7e97cf7426f72fd48ec7b59023ba9f11537d62d69d1b7b725ce01f480fb38b7c642d7c43f5bcfca6a19545739b879ddfd2e62cd0bd6d5af2aa7b0c1ee6f6925e2d44173216231d3e2c3a2a6cafd0dfdbbb96936cb388ea286829c431e85d49dd68bea82cae04ee4e68278d590f63e36c2993eef994aa95426d1afc26bcdb9174303ed2b08e4797e95d5ce81bed33acca051bfbcd06bb073ac97da446f1c186be926af222792210835e689bc423e3afbe1728b96fe5545e466bdc0973ccc69d1b6c829057193a097e1a7e8bf326857442de4a950d04c1359953d8039615c22b25102ca8bfbc3491fe137f1d780aaf61871ff7d28ca42f7c2e2e74517261287ed0b749854d310289d2ba4995b848eb479e512690fe4b34192698f8a93ee944006c033abcc6c775fda975a8277276b41315b7fa59d06a460fe1a42b36aeb94909db18fc73695b3236b42bc2a532d304cb4a8f6601fedbec30d2bb4d4bdf5f19547f84b25d29897ecf334461391c14ec29133c93f0f407206bc2cfe3dbcaa3f5abde8ba402a472cb01e46a63892cc40c468be65c575e62f0970d37f6ec1b865ca36a55115410f4a3328cd14bba9581a7a4d1444dfc3f5bb1fad28cdf5d4c96994a620e0941be6f88dbc771b40b7101e9a6d61cb832a21f225e0a9f33ea474d0bb2f95da999d5f86975d9efbf5d3b3887890b5a135a8720bfcf23a7dc52aff3bb4494ba41108302d5a34f93fb9ea7e7a9947996f90f296b41736d26ca1e9469d9399263c87f81216a40ef0277bb59899495b30360e07ab652c5e50bd9949aa87f1e3dd20145321994940de777bd1fa1961fd4829bb5ab538a20d57488818d217e521f89b5be0b8e6da5f4441a0cda3b4eeb85fd979ee3bb9ce365369fcc54b6b76cc22c9979d0738c04e1fdc8b32499b3dff7e1d194eeed0726b1fae1c7f9bec23184bbf6988b323fa20dd804a0d2b18bb25c7c58d0f828065dceae3057638413591069281c92837b5a6c9c58e475796253d7beca3d55a6f5bdb7156738129a02e1c287c6c261ea36f87049384859dbff7aa44f5ddd71c8131e6890188c6521a938914bb12adb0783537dacce760c5816f13cc80a00f75c0bdb86fab67591500c4d41be4395ca2f4784c522242b8b43275a9fd53ec846411e9799dbc72fbbcabfe30aa459aab6891d34289567595f49d72af23f58ad5cdd555144991056ecaf3526050e731e2f678f32c9679d7ea48edcc2ad748edb1b9c2287444a762621404ccd37ec8a11d598733f2a3c13795b9ada5601f796b02fde8a25fcbb4530ea88ef6940ea19d230a98125b6d77a1e7a709395e92a3d3f2a46c0341847a10a2f20f410c79c0b10948d2edecf18df21e0b16e18a6d55f7762862691a9d5eb2c54759444241375df9240a3f432c9528cd578ae27f715b99f26f2f180f435ee3d5f58275fd45386a5f963b1e7833820950c058dca9715eeb857d492ed72fc74cf82c70cba990acbd28e598b818dd28b2c99471576b5fe00f32936ff46e8f91da87036a7c9a2f0b9056b93a0dd21db69366aa2567e313dcce3d79318aab62c8750b0af5f7ec271d269678e55f188d6eee97ce8d37cfe01cc35720818a8b43ba6b06ecd413cc00c48784eb13ed6bb1d76b0bcf5c3b92efe940f12ba1e798211b83ffb7395e730609edd322e6aeb7f2e5106ba02fe68d9bfd1418c50f97b203e9070ef034d92b3acd4e9462a99c18d0ee640fe9a4c41e411679946c881b3f20845ec4d7dfbf4d4e27ced3afc7c71086e219c997bf86a56472bae2725f4f397070276cc1c043c10db233c2892359c46bb6be7f7c477fe98a803241abb5c0c5fb1269e9d71040f76f4b6b482b7341ef11a174030f'},
		HypertreeTest{'9f86d081884c7d659a2feaa0c55ad015a3bf4f1b2b0b822cd15d6c15b0f00a08', 'ffffffffffffffffffffffffffffffff', '00000000000000000000000000000000', 'd0ae6456d27c8eb3f2bc8a92c5ac678b', 0, 0, 0, 0, 'bdb07bb7c73d3641b3add3843dd34b6ee2f740ffb715414b308aad09c7dfbe01c4c98fc7deef92ce0827b0df3ae490c8454b6eaef357a1016e09cb8112d9e221f6b5cb271fb9060629653c0057233edd059d0b9035697aa4e2abc08c5c3001529d2cf39965d7ccffde2b174059659ee2c025ffe931e4842753f47db60ab6f377c072ae6f6859bf39f1408623609ee848b15cbb6ddb66a3576770f23ec7793e140361166a848cb3acde88aa22968db631229ac7e807c641e6241c121da0373abe5dc6116d71632b2f82ac238eeab0c4c3162ce502a62dbd7c0147e81523af3376cce3890a075918a2d8996ca7cc5cf8a3f5d0793b3e47f7395abfba7552dcbf66697127ba45b9ee9cc0d652d719d615ac699aef2127dbc0cd464590120f4e1d01db5bb640dd8a7f63e1d700342d103a3e54d84abc28ba43a082818ff0623acc05d0299c37b6bacfe1f613f94d596abbce4342ec2c5be0802bd556e9718503a1cfb8f4f602757852369dcdc00cc3394f09b4e23d9a371f63c16d0e7f8dd84d970dfdd2d27163259c9d6b9464a13abb5ee73ef1e1e17959d566f1d98121774318bfa40b8c035ab7a0aa2f6136a5c99236e479cb9fcc1cfe2335ea1cc322dfdacad2446770d211856ba293b78cd707aaad890f53dda6c1ffcfab64eedc4ab1746afc6a74fa0f45e9a9600dcf703ec974804c24a677baeaf7772c704e755c48223f7c942a9d677cf56fc6fb9017743a87aaafdca15eb1d78114ff8c2329dd67d6ac0e3d7bf5ffff45910a1fa4831522d18a7943d6413819a4fa14e357bf8c09ad51bf63762cc3d184a2669fcab0df2af504381bd3a5e6ce0509a1e01d046030ce7b742cd06ab122b60fd792c8877e7323498ecee0ea0f35022af6b44f805b48f1fd6a1fc0366d09d8f209de764556ebf2768ff518a0078bee9bb4ea29de8b86d715598089e3eb1a6bc8986212b6e9f707019da313f022b4dc78dcb29898f4b305eb2c98dcee4a3fbc3fff8c469514e6d2143b47425d4d95f7f7ec70138a863d60508c4bee6e228fddced410c72ba5b5fccc0939d49edf6df86deafe450200a7d9f7a6bcabb26436f8dd9670538425e45e8badde25d32d216341a99609c907a464969d72b253172f52944e3f3c436cbd70954f1281711478d90684aa735a968dfd044d0f9f0705a281db960e63b9d0fd6e460824c68628b1ce4bfe8d3e642404e8d65196eecca11435b0a31f1963d796fb08151a669d54ed62a0c9b4a451e6c23cba5ceaa4c60185221254302c5b193edd9be343518aafb63deb950d01f4eeeaad5e5fb7d96fe53e5cb4d51307f90594a11ccce5107d623270e004b56da8f62556f50518526594fbc4ec7a08ca2f1313a91d53e6735db73d38d809033f1e19501a4dd86891eed172d50b7fb02701b0fe98de374e887b34f74a587f40fc2fc265f6874bcbf2487cf1fe5aee36f3f08996450f848d1cc2e0c44793dd717f55866ef7c6c69dea32b61b44daa99f5c435a9834dd0422a6db37bb54f0b30c224a83bb0c059a82a2889e16542b4fc85e0b21cb53f295f40f27ce6c612b477da6e25670df1b960ef5385e59521a460a14b9d6a7590586eb5fcd66ee7c98cc2e34f59ce1cc8725b981a6c0dfb203af7e7de9517e9c84314648f57612c13387e567b626cc8537515241fa3ec0acbb6053986adc8bf0a0e49c866b96f9c5933b82feb396958cff05c8016a2749882fa464ed72726190e8796b4ff5efcae2c4fe2dc6b4fb36d7a77f546ad357cbdd88903f6cfae8b2f0cc330fbeca4d25716125527f08fad7bfb117f682a188d68951899a94efb568a7bea24d28c06a1f0ceae4b2500adecae3d6232d215f90f55318c4df29e964c7aa1da40a954693d6f6ff3224209bbdd23c1cbe73299e9f8fc39e5251e61a0d38f0638253e8d8f6105c746be5207efc051dfc08bce9e8f03ec5dc7a865ba88ea9d1368f00dd205283866ed4d0e63e0544104b64c195efd2ae8fe5d71af7b07e00f8455539d8459473a6a4fae119d470ecb4eb7ea1ec55a6f883c6e5001c1c37fcea6411d997df68345cc44c44516e02b936b3d0721cf8312195694bf6b098bf8450cc838819533ff48774817910a725b0f56c52472890982e114eeac1ece08c7ed72c4ab1cbd35a6b1aa0d4f152f33ed009744ee4c3c4efe210ef78c7b4e403a69ee03504050a8ea830ba11acf4692b4b34e04d223a18b923e0c19cd3fd2db37cdb5b31c09da81a0e6772db083d8846c5821c2ef2174d0e0b51c4ff4c66aa9ff49d3d13c5ca4d2523ac877c15398aa662c4b91a88c4e69f0eff0e89799e92964a71c39258401789f7551f769fa8e2c643d96f6fc9085a817cb5ca132e3a949b2471c984bcea0914e92491d4843298542f57ebd0c1bb78d9162759a23678ac5bd638ad9d4ff0eb4cfc3e67ea6e3c014a102916e5e7902685ab54bba67340c8e51e504382a00910013d1cbbb5aacb628ac4a80f16e3ddb1a3231b78fa19023da5b53836aca60139c4c350fd6b0c2bdcffab67268ca4891aa4f40a84f750e4978061323c5e059b225b4d67aecf488e57f77fc2c42c3fbf9bec2ed10b0f9056a3278fa2d96aa837e3369a205af64ab340db37ad8f1d2c2167da0f09275e5508da7e8eb329e1d364e1d105aa0885d43fcf1e7dcec715d4317b331cf669a3939275291ea910ebc37d8597c3b2b3c19a654839002f8e007ecbfbb4907418d30535adf78387681eaf94a68a9763e697bbce2727eaccc3df6f3df68e91b827d2190ace56f207af3cb3f18e6ccf43e273e0d33582fc1e8ce5a9f7b3051e0794391403ded1562bad879ff3637a9718e46df0ec5e00e1e4551ab9d69625c14f9f20cc3b735805ab13bf631be4b274664e4ed8cef75db25682901190e369c2e5bb95078a2a5cb1b5e3fce0081dce6a1049b57711cbb8b94f471de53387d6bdf849645d2ad489f66d9f5cb598e385e5b6cb026b89642e01101997eafca4c37a722f825add05ce55f91b1552e6332f521a8cc7977bf9a9758e776f3d65b519829888150c31a7b74c5ea7f1deda4a03d39f918fceee0677403b9c6f4c88a9c499c9fadb56adb14bb773e1333b0d55043fbdfe91234b90d65d8aee11091c0b445d7869ba472716f89e38923918736d824d0a39500ce8cab62d12ed09c2278389cc41ec3def980f15cb1198361a25c4f0b6a637695354e3e0793bf22b758f5ecf966fc6a57fd1b7bbc53400cc7268a3455f34b8fb45c1969964a1322e4227f8c54ac509b338355b6652262ac1bd545285488b33affce78139be8ee10424ea82ffff96ca6eb511b9c854fe8fa73aefc89e702fac85975f90339654d108f93455f61ae1a23e007ae916b399df2b37206ae26a53f8f68f7b5399cc560f93b0d348f398de02d1499f0bd029428034e477465fa600c0a325f2386189c22f711c9a80e700d59b3f2d7cbddfa50afb5a41c16db6cae77dc4a4bae22cc22b93874765443b79d5d89e8e9ccd50d2e9cf4eea8313d1e64b55a6b5097f45372d05696713cf0fb84fa1988b100645430fb8485b6b52562a601faccd528dc22283f788414b78874e69d3f378d49d5473cbcda360383b33d28e2dff21817f33af8507e60c4e132f9b92a8b5d1d198711c8a65d3b34252eac3d92008b43e7ac79b382ce6950b8e7952c0e59744d4de89550cf272392134bbe89995066a07848aa7eec66ce304d19cda806352ab5814a2dcea47085f3553de41b546f1b3c9c0accc06409616366643106b0433a62d50f5cf7eac86f6020f366a6a3721e600459d0ca51eeed4282c45710f47486f4f5c404916a860136df7a3abf6b298d112bc65563343fc4695575615580147e9b66f4b0203e20e8439d08f2230b48dd0b2df91f9017c1d0fa2b5609cfded8212c2f805aaf5a091476a8cdf385363f1e02e50ead5cad01e019a6f26873e000157d14c974e756046e3c5dbe2836757469d0356bfdc7bd11b08dc0b72b040abca7500fe2462cf164bd3b264923a1d7ddf54836b0fa32ed53c9efff7dd87882ebfcfab63a2e5eae0e36571afd6d74c9ad034e436db0d20776f791fc41a78621d4626458e1f1789f7d1fdadd81ca1f79682be45ff6685e66bbc092ff91a691f1eec12aad04224de2af968e96673928cc091ce25898d6198d9e82084d49ac03fdf5db875dc5b90a3479745e12c8fac4d42c9f9d65913f033295d9d75f9a0f3213af70ec7cbaaf56d03ea82a9fbf70b845af52a55fe736f8653e90f1cd5a0415750568cefc26d30542cca8fcd6c4572d702ef023d294df100557792057b84172cbf17b71a55cc3e399ceb66924a78927fd8beb6327d099774ea022af5cbb4ce8920b92b6ab40ae49eec27919c9a712bd7c91ef31ef069b45887bfffac54f58b1485afadbdc17e246cd3f39ed0ca9e87214eda261543c6b6ca8c7908118dd883dba5eb82d55601723addc8749b7e2f0ff7eeae116d8beae3a9d19f79df5142b0e71444d89be0c6810b2f874a1e7d0683b6bdf69f3b4d888bc15fa9551187cbd6905bd005def1337b7658fd6835b6839a5bc2fa13a4d0c740f669d598bde0a529029d7481a8d65faae84eb3af2ea41ca2c42b361d728029be8be1bb9323c1905b71e7f7b2b4de998de01cca64f7065143c1c8271f1b050c1875f40b2dbc227e29cb3eebde568b92ab02abc07d6fb464c1eb85c21624dc1e13b64465164103fa5827b03acfc967d7d8bd683d372373b42af8bb559b54c320cb7468938881630572a3b55b0d2d9dff27ab2f4a237c731d04b19af163411ed1d274776429290e0c8da3ff7c9305cfda1e129b9938b4214a7c69be7ea86b68c7e952195f665d1329835791c05e55e5504711d27a86bb4e3ffa82989d80ae2695d0cc705bd1e0326b773cda54ba1367447b76cb29706d70aa46990ce25252eacab1dc03708301417f8842dc7f3c3821719c357b921a7af02d939701c8fbd8b2273e32f0c58ad77a647911e65d2c4fa7da072426340b9f3ba1c7715d78f2e79de29905fac7ea41fec2c5b30a884d90e582d0141ad5e841767eee7d3267dcf7fa269609238e9fa1702170ca17e50530e244f25102e66604f92d2b0b9ed97b1a2ee31decc9617c14b60fa557b020bf02a31bfa1a1a1d2ea2f522ef297c086104e6228c20f2f0630647a533802b187cd3dbe90ef2197c9b27782a24ca9b3ddc8804e40d16e8fe1fa4db5d601accdd65e1c1fb4ced86fdac6afcd82b66d3981df611a621e70c238a98e9402e69fbbc400b84b20f03f95c1360ad9a135a009d6b7e1562bc35af9706cd253079468b03de99727118db5d5cb6843a6d4e2c2a62a8c563a82be6b803979da611070d1a759e07465e92d7f019e8df64f755b43d6dcdadcd858fa8b60a1cb79a1c26f14661f884c3fad59b33873354fb940c13ba1472f190bf29355b8f1094dba98d7f1f5cdcd0da7e03629bcebfb0cad5b9e62173a272d5058d3e191923adbe55f1d019121142d5c993d3c24ef25c9611ee716584a9d10acc66b1d10b82a0e303d85b376cad25291bed30f244eb9323ea0a9ab0e5481a5fe0e3979d286f472d407603fe6fee40b541d08bf55b7983811591f26832857972cbe170aa25f725f8bfcf5ef80f2e713c13c0bebf2b6892c9c589c2fc44404c3283d68b2fc36e469bd9e6ae3f7994f8dba9629a1c2b5c3c75e4e79ad988b43375b26c240342e235ac42ab2c26d8b5030425972c5b528480e5d13a0693b669c57517c1d1f224ebdc0218dc2e22a73ed71bbe14725e4d004ea130443920d1ac4bd08d56420d82643b2b70fa67db994e314d2b581d9f050ff1e9289b6a896b210cc0a70a352df3941b1ff1a06280de5bf4c1abe4c646ada7dce96bd21a0776dfed803a2648fea77e11e7dbf94143361a99fa46b4cc93ed1d63b7bd8a106e227e8f174c60bbf76af26aadaf88e2f3512d05151bfbfa375fc92a82c7f62ebf2193000c37ae6bd10418b2d3f447a667231c8e65fde7bc7c0af84e5755c9546b9fb7ed723be9edc20279fe029ee1d33560df0cf7051259ecf274ffa794b97b0d3139504cfdbb40c6ab803a9900eafa9e703b69829e28dd4382e90db8d78cdc0c1a2aae049f2c2ff95fb097bfc5420e8c7cd3ba07d8ca18c9998546aa1c7bed4971a51c46238c9d8f37bc722a3f0a9729bb3cb24e2537181f946549a41cd9617a640c80ee8fc5aeaa1d3802dbac9430ddb9f2b6dce1217c28128799e1e6a52098dec1bfec95479ca43f07adb978b0daf061f342f076871eab64acde993ca82965f2f0bcc0d2adac23e17326d0e18701d5dcb780213fb0dbabe29ba879f00e012c8faa441732c5c20ef529afe05cffe84471de6977497685f6fd1ccc5155e0318fea9a53df877e2effc37a839154d6da70c8c9abaa620c2c97d1a88b4f47ebad6a5be7b277922d1a1fd2b2d825df19562ab91197e98d9ad90a4df2bad2a089f23ec2109784bdae8179aad1f2640561c07602e1f58aa778c26bff9bfa4685a67ebef547c3a0b94879d80d91db1825ab3cab7a3d55f97e0e36e87771082b22d00c9c2ef2a34e1ea54d27741b0c0b0ada17fbfb725cc04e1f56d4dbb4b44731bf53e078ba33a03255141072d392502761cbc344579d595cc788387e016267ccf01714b50c6f237d3276d26fa6398724028d8b78207fac8f89557d0c1ada0b6ee769f7a7a5e38402ab65b07b1b74b18f380437f2cf67647795d1464705bd7da2b934a333908b880fd6c3ea1923dc7ca19aaa4098b1b51193fedab5f3ee9ab425403b6f96e5272a2db8fd89138d9e5b5f986b4b527a2c6295b8daf7c882ea6c73e9b63116068a868ea9835d9ad78011033abe34c7c4c6704c4079f691a5ab6d9bea59af1715b7dda3e297104cc450d5600b1f084b71a751f6192c71e25a069ead548c8a00fe0b87833e381bd2babb8ef1f8de17a1cc19831692452b577f6b57e263d6b994b0a767c4c8b5ca6b3e1192c8ee9c2bcbd21a1029db666ec1f4f4a611546232d9f73eb48a25fbaa8673a524ec86767a8cd7c462ac70b0fc3041e1a9630a43f978f3c2a957df32d1b304aa0245cb81b117d9b3074463c553f208cfc9b7459eede2c099924afe35a68315573eff819cb680a8369ccaa994ed9398598425cc5fac6174ac3c224826a27668bea4df095ceba7884bbdcd0da250ba74eef06ebbaad0ec2ee52702a186042da5d703d5e2b1b25b68f66a7479b416b215e66c6bd20bfd874a478418ac1ad1d48862c5c843821992b1fb071fb70e6b9b0418540f935560706b51285510a35b73f8e838f4dc7f62cfc2e0d06c0a4d4f93149b66e9775891c98eccaf9a52ca502e8e19244289593d82fac8b6d4bad1f5c1fc6406b2e545ce063077005977cb4fdb2fb505faead7f70da40e62a38db57a692131c4052dac2e5f176d79bcfcbabc77123e86e083af62072b051126514a86179ce9dd120014963d1aeb0d3175f886ab7c28f33e340aea35fd051e241e57b58445e36682f4286716d0f05d753308b417c26e18d7320a4de2fc2fa4dd7774eff6e19d880af9f8a9ed7b4feb844f1afe7937683af50b3a61aaf143156a7a835595699cb0a349290def8af1c66bdb3fa9f60fce44da85fef8d1b6c0bce5473db7d48707998152fe575813de2979c2433cd365b7ebee164ad34691b056397c1d1b7873bc05e8519d1277a481155a6285e6a78a0480c7946d22173d2b6826b196509a126c626895f476ba6d75313e52683e135bc658a031992ed79570cd0295617c7ebf698eb18682975e117be5854c825c084715c20b04bf8f155c039d156fddcac189a410a81d7d67c82e4d2b25786d1c70949858903e1e484a13eed5f8e9b5e9335885deebe999a65b92d72f036bc097a597233fe92f350f53badd59e54f044a7ee0823a28be79e2f408de25bce972e6ca65d267bcb6421d926567b96ff23df7f873b18eea37515d52cf371c351cc97f30646aa32c3fee766bb812a75f1d3c0763a9a870558855b7151fbf001b323d855f84a4a5b861ce5379a91443316499dd88e2becf38d9f5d5332c5ffd0ad901ee2b4b96716821a780833ca9fd083fe8a959d94a1528942d473f44f546861b94763a59ed767116823b8145572f67f1131c4c3cd79f2451cdca2a4b0cab7b67b63e3e95fc7b59e60a9c519ce2c125e12889610db69c6cc892ba71cbaccce3a957cb5616350832ffd34f32950a372f2e729b6a36d7e05de4d901689a6aa7ec23aac7dc7871f10da9ffe5fd302f358b38a1a0752df3e26d4498253aa3ee022ba1f5ac72dd0ce34448d84408cf2330ab2768a70c70a27edad55fc7826af542fa9c03d628dcd033f9259fc69565cd1136259747334e89963ce400964fe74bf344c910a9f75677a4bda89d1cc68c68ffb803bbe391076d84a5106b19fac5ce36d68cf2234114ebb322a1d0e87283e95bb55469cc7699f45f420993caac654b0310ecacbd560eceb72693747756344d4c4c311e42edd70947787bc91555935bf566b19bf2c6189b4346084c748fe708f963d0b5cb0a3918562c1796365398350e71e200c8c3d701bd6aad557a536d6ef9372bca1aee9c02e50d920f7f7a00e971dab02c193e321e927f3605e340c88d8e7208b5d3a4849222ef9c15ae3650c579f636eb77913c78cd58c3e1a7aa06d796e8c46f9962fed835e09084d017d1440c2f8108dd89480184e2740ec7f1003938bdc80f78f10dfa7452327e2f74c1a3f57be1c1572e6558708183c699053b19725f1506fc441d327c26840af7780f48964bf77c9f7cbddfb78e4387a636bcef3e03f9668c92bc56f09b1af2db9b51fff373042f39e5ac3da77cdd53899d04a0e45daec2d32885c42a8bc01464aa478eb3b7801834689ad1fcf29ec1d645760b2661f37f4df41b4286b32b48251d8cf006747e983a864377e357c5dec54aec0b0cb8e9d56260d53a96a2505b26d1ff2367ef5df97705f4b8a0d8ef6bb30361d609eb289c21f0db94c9a80b714675435d1cb41d8c37c9bc271cdefbc67378d7adea47bad02b7055e9bb3ea1e851d17f9ccf5f931d67ae54c0b2d61d7fb87ff046f431190ccc14b3aab18dce1ca8d3a4b34a5406f644770e846e5f3fbb0301ca0b24b90d972c08a8e328aac10692abd26c557307e51f31512f6d43250767b12bbf0c9c5e4aa283f787bde43908b2493d76d8c808054bfaf5c3e190a60701540f936f9f38d4d9b3dcfa5191c2f8e95303593fda45b7fb519d466d2084baaab06733109c1b1a7d347956e7d4e6a0bcf4261c0f56bf06f6e59b92b7ed02885a8e93b1ae55c7bc0e09c7d3580447ebddb75cd74a88d77460ada94e46c54dab4a278c80a2d12ec2408c6ff7471e82b9c435123ac484be7f0ae2bbfb82260d96c1f94a1ac6dd662df68f82ac5fa7e1d715b46298026f1302d11302cde971b2a7dfceaacb3538de1988eac8f2233fafe184260b3747e5adff450af1d73be0f97e9c4423140de37e93289b7b9eaef4e61ca11b329950a3b5719ccf4d24784e6090e7d418886b2fb30093a18ca88d39dd95d88f1d24930c9f6e4d50cf7daf86fabaf197835e1367d9769c167187730c4d9c5ca1a123a6dbf7ce1506f16c0bfefe582f6a3f6a41cb6e7e3ee182d72aa4f00fce9767e054b84b9801854ebb1763bf6fa5817a8abb837a4020c254c341c26443e9c54188b27e7d5b72e9dc588de8a7b61357f95a41c7dbf7bbd9485b5630717fb054be9797027ae7e63beac2eed34978d489c3ea2383702b89d8beaae4c192385ca865be8d3a9bd116410e300edb57ab8ffbf08ae68ab5a3e2289f77b1174762bdffcb43e0716c035381f2212bf85ceaab98c4717d36061216f1c208be3d902b408b32d3ed099eb048ce7ced603778b3eeba3e751fa861505a22f74a10011eefbeabdb33795244690327d3a96fd079dad0c2c8b0c7e8859d76ff0a8f28b9938365e85b5f02c8ec4a45930699f49a7d0c1d8f966f6f446c598933ec3fcaf8c87dc2ebd04d703105d972b00bda4317bcb5362b583b362916b151d09cd50d7c8eb30b4fc5c1acac7c340df85ff436341dab1e61b4d002dc06637c5cc06b5705c06e58593587999cfd709cc25d1736b3786270c6a26f75640b354c345b1ab71692cc37a3cf1e9172c5d5398dbdf53cd4495b436e45b4aaa8a520d94baa61e2016476250264ee3a2df82e73b6aed4065446804f717cba85c9aec808ed8982bb1a204e225ac5649195a45b5696c59f7b4e00b3e5f88491e8a60d748a6dea81cbc63055dda3ec6b58628f7c6a650e1f74e3fb13bfa5ff4f7e9f5fc61b7a9d83a5ee38366957a475b72f83dbc47d34cff119f7279665ba15c7aa47100703a6e54d2fc2b284c8707e50e4869a1da4098363d8658ad78bd8ce6ea0ed6d3882c2ae5431e1e74233d84c418059d5daa6ab6edddd7ca1ee9f5279ad23057838669e50a321cd9049072879f3f3f3d7bfc1c65584b4ab793ad69bb95c05d3c3e491ad7167b2c0815c6ded5c70c1214f95c2e7c876812c7f631e1bfa0fd76f485b74c4b657239a2a5c52fe28af1ff0d7171d6f82f34060ece3d604615bbc2d9f7dc58910c0aa04e38a3b9abe654b60b48f52cb90c3dbf2386b819f920e0fcb0fac382ab636f2d4a22e391585aef49c99723d7566ec7733da771b5ca74483bbec0fec7f843a943673280b05c3f604b307548d14c88ef9b7ae2ff6072b1ea68f9de99e88f834c3686438c7be74976835eb3e6c5140f65057b53b37bcf1c869a87973b325e6457280334cc11fd7152e03b5c7fe8662c4ffca429187cd287d2bc98a8dfb2f9acb062ca6770e7846f13e528218e4e55a46e4615958ab672fec4653d9a0d66ad7bcae8d97532bc300241ff3ee32717a2303df9d2471f34bd13d647ea130742d688dbaa884d604b9315dcf863c1fc8d1b970263f990cfe1cc6633d57f9c15304716916e62d126ec398a80e1d89d4ae535cfe60f804b31f16feca8259f1149d57cd9fecf2056b5497072a77fc54be149b3c7e17dad77c1b076c8350ee0f9ae12bc887248aa109db68dfa7e970387c97c1d9a2488ff8c709c81fbcbd54f8e656e29a1ae432b137a02e95b9ff75b6f46377b2c4d605317479cfcb88a1571af98d3daa72683b4534ff79531b8e0361cb658883500d0d6cfe7339c687859e78c76940539db432845229dabc3ac40bea4ccc8119f8409dcca9bc8669968ff80a70704782928cd9628843087786e45aa065479064cc8aa259fab45c62a89e4f9b9a6db40812796be2c9282ca7a3e803697f60da737a7f07a0c959b1bb6859172d841c6543f6d4affac61401bfb9cda08219ebabc925d895b4e3070b5d37fcd2f7f4f27f05a6dc6e8b4a1221e5401b7647fefef41b8c3d82bfc2f50c55cac4b0bdd35fbb47374c4c3cea4ed7a3d61ac17eefd1978604b199527c81895d2dc553d9351383061daea78fbd750886bc04519c16f35ffd2db9afb517ae243ede95464f654602ff477a675cdeea23a802afa5d833a331efdff81873fe7a580b2d3c4e4efbf7bf337ff4bbef30519ee13767956f958f26c31be3e07064dcc24dc828acb2b3815ae18239d20bef11853e0521c60aa593b3beaa353c86701137b1f12a4108c0804557a825cba2426550d516e6e6a6e2306cc61b2677ccee45bb6a2968cd7652527f036a8e969391a9eff2e1c1b9ca107bba84af276aa4725b2f9f52e072000a74654ed7ba65cb048609c84cb4aa5e24a628d55b2da0820655b916b41c0e1b6ae6736a6b5191da5e6f2a82e88f39f2c598a89ed49bcd39797a0174214f347a76d21e30094023c5d0ac778b77bafad6ce63d38f68f4a6fc9d33cb029bc5e40bf0feaf04a3b4c230fc11f10700464ad35dd82a8aaa2acb6ead546c8028714c9979d189abb4389cedac878c05fdfc2dfd0a37469f4d2bb7016c2ee136fe1d9619d76b4f48e063fef6e9e9378c255ab2ff52fc60fde2cf88c91decbe8cf25a2e58af99523263e843872a6d8757d32ffcf9da527a4a113d2408b14b08dcfd8f5d16e9e620bff6066e0eee50dc53d8f56bc84f9157efd2a5c8a45c3d3a69337308da0471a39cda79e3a3bd58cd5f0676bb0e1affeecdee449de62fcd2fddbb9f11642588cb6701e02fced94e5a839d46f1966ba580bea066cf1ebc70f27a40010ae903c6b8b18ca10a7d9e3b90a085b7f9debe74e8b440894c20c0efd48ef59093c5c730dbe000b9992fad3881b067f424e06a43f65002099efe232a37bd1bf91d81f1a15e0c90e43fb92f2e0496922eb6e42df71d856ecf7898ada46d5cef4f4f732a794c931a67e7459ac12a6d2fd2159f9822a413ce123f5aec4324ac67acf794bdd27b4476f281114bad247712f3622bfeb127900bcb1eb39566329354196981692c5461dfb97d097f3803bc69c723776703cd54eb814d1a16cfac0c099bc774c289573001eaefa7816bef1e5fa578b7ed3603e73c6db2d41629959bcbd2e6a0973155f32ceffdca1a42e12e44338129990dad19e79d0c39ede92dc6632916491d9ca880e226a30ac53f957fa49ed7fab84e6cf62adfc3e7e9317c42b14748d8bc4bb6de3a162e60b9ff3329cbab1606c5978a2ec016ea01b2977191e4021998eb3aa2b87a1fa5ef0af7da3e608b6e57381782e1d2792d1448912d79f0e3b8298d9d00ced9b32e592a4f96562d8720b9d2a49840ec676a067f89a0c14b334e7ce2e967baff98cff375f1e76844f30d9515a9f0336cd1c4f37f686da7c1a2a81e296d89446f0eeb4e95122de21175a815f6c6f1078137f120b47699ea1ea466e372220a3cd57ac514c84b3838d9f0a9975a01da1a2682ea9d3ec0c5c91203d933423315c0b73cd4ffdcec90a7c22a244342554bd99d545c8d5344541e654beed4414d7fff0707d0ebb488af6f55bc08cbb56ca491b732ccce2dddd6f39af7be52fd5bfc451248d3122094f86fed479f186e048a211791c6a5860ee9d28165463b5927ca03b4b74905dff01243c5404a98140748f6d1dd85dc996fdb2ee0949a80d5bec1294c6aeabaf59e3f3860d2a4d5a4595ad6684608d7eb946c63b65c187c561291e1013b472ec862ee4e1413255eb8c68aa465fb23365d96e10ddd4374829d78f78d6aa9563e75e15fc77770b2c6615b363912c84b862c0a20c2cf5c7f52b78edbe7a5ffba85359762c28c47a1347a481015d5c190f07184877a2d4f536ec23dff879301653247d48830fc3003f1bf82fd0e90d913fbab97079dc4343ce2a423d92d6a9bdedbbccff060f9a7e2c7ccf06cafacd51eecece49d2e5fb69cbb678b28d7a38f8224554f5eb927bdce06ce152c7b802f44d94d82ecc97972a3a7e93e9a40f989e89e34e845af4d7c887c42a836a2e458018b1fe1c4bcfa912ad708222829105af05c689aa1207178c4838f86941aaf624131c35718e8ab93720092324bf87c4baa0ac9f9f9b31aff3556b92acf30545bdd78ea402953b2f48280b4a6e4554279f562bd7de609689b3e199e27187cc9d62e7b0a9280748d5df6e3c1036d6de0b0008b96387949d92e1d1cfb25058e52460456a26ddcc8f28e144c389e1cecc6ddcc9cadc9354887a70a353859b709dfbe29d825574d2a21d8c3406f67768c846d3dd67442d7efe921ffc8ddaf8a9aa0e83239978d8231aaa86b275c873d56f95f3b9c3ae7421436df242b91200c600169b8438a6d67ea33588e8a384437b2750b731e34deec1f73db337080c6d96a69f1dbc45b8a6ed663223ccf2b0aa869ae478260cdd5f877948034569044d4b6521f843e85cb5be304bd8be764a9b553c34b7fa7584a1fb1209e824e42a8be2216e49518654e8bd8f34b5f80053a8af17c804e5b215520e81fc103ec657c90547a109fa6bb318b49830949ddcdde94457388d880441f56f0641ac3489870606d2ddfb7f327158c8d98a7296e53131c89439d8c6902d6341e55f799b2e42ac8b7020b68654f63e5578af7e97d63c74ef3ee76c11b6789e4aba423cc177bf97ba10ff3bf9bf2d1214bf758a4e1555c4fca811a1f8da4e3f4484cabaf44c225856d83d06a7de9ac78ccd18510809b4f6ffc2c8635b56a2f6c45051c1e18f4ac072bf7ddb5812c33efaa475e191965fe0fd4e1ed42e67a182fd99e709750b3e209deae34dca3f17027d21f24bc076375f4524c2cc1234c3151f94de8fbe01ba78d5b39e91d63ec6ecc2b9e8e7ccbc09390afd070b62da682962e0a60c00be533e90d234eb26d1ab4b018b521666c3ad4c0de8a32ec953056e16b17378a56363dac41902c49220679eb15856ebaf5d7daa766683a25760bd69a51b92784339a3bae16fef520c7232b65c2b1b2d4c641e2dc748ea9e6658d80530fb00d04b49a585506396461ebf0ff19a1c495dfd12a88d3e7d5f104db04d8d3b41c6253c5bf06dbebcdfe5557e62f98483b72ce1aaf49a8d1e6ebf997dea26445604baf0c660f6e5f3b22cec154fc141ffcb0fe49503cef70beb4658ab6e78cd0b8b0bb0ec2ed42d6ee93b6d23006e618192182813cae7fc94e469cf73fa50a3c230e7aaae172651070654a98066bb08f7159e64d880dc261bb6772995f1fd23d78823bc73cc7650703c5b677c1f8e0240227de5712450e0b6d97454a99870eec89e5cce5ab3f024f85af751aa132dbdd9db1af5052ee25859ba23bde838ad19debbb45b2cd397629d567ed9f6a10a219cb02f6c153451e93caf6caa951200afe410a95ade425bb67c5bb0dcc32e496ed92292fc70bab055a51c5213f0c529b32d6b7c3fa6b9c9ec656e3a44ea928dfa1c18d3e5a441f06c43d298ed0588899ad6b012d907db1f879244ea3823c8e30b6514ce6a849fd2dc9a42a5d480a41ae01babbf227341f3cd198e93775d78a97a5880a099aea902491f19de3ecc993ad5a1e73f8ed097ad4bf784c9481ff28a233ce678f1df412106edd9f3a336f5806e7588fb75e397388ace09307d8d2270d9659ec1b5dea6ac48dcb2ef74949bcfaed36096753720294c5d2d93cee19f7e2403bc6517b2694df205fce1bcdb1c24454b97c734f6c3def54b64fc528e546a590c827329daf9ac5b8bd5b0cd33aed68fc962d2c5db360f85842a18c1585b457455045f7e508f0da17a30e9fb18bf509a7785a8924d89f5f821d58608f2c6b33cb2288edc8dc0dd08b04c9f9348d9873a2766b98345430ec7d1ed1eb645141ece57bdfda2927ba937b1dab3ae9b36d1fa5c314b43878cc7025cb65877b373b7fff7a1e5175dbc1c946989c790597b4776a01e2f6130f26f8ce1ca6f07f21889a5d23855701685f45391b30d11afee14207d4471d392a93ea3d0b58ce4364077d2230199d7bb14dc2e8d0f688589ecc9f6a52dce0f86f23865eaa6dd1afae32da9ae43aa72db322b40c75c62f0296bc7264359e9110337d0e2c9bb4322a86c0bb97355b08678310d32cff3541ab492c7be269240fe24cd43cdf031fd696e318ea55a2e3c55c74c773f7d2231fcae6cc0e9a5ec44464681d6c8f2d0a5a2c23104ae8214b8c6ff9727ec9cdbce10220968c3538afbea1aa54cd89c113210a52d81ddf2bdd706f6ead8bcba605b15e02f738699cdbcfea927e67f77f03cc1ff6f22fc6a373a1833c8c4f75620bd2f33a880187f113fd3634f30819a13d0ae8352ffbb7fe4ceddb08f50302b43ad89ce916715ab063ffea3f235b91d39d397d26be72d20ae7f33a5f06ceb7b5ac016e004690d141641c23d9d3eb77573658a53b2d9b21a3cab13a63a4fa2edc1697a831f8bb53aa9597131bcfdbe1073403c32ee2a0b671dc3472a577ebdba3a9eefe9158ab2baf544dbc5d38078ceff13bd19ba2042c8c77cdf55f2fe0393692f1a314617075289ca48b3d047959084227dfb58522f8c240d8ffca50fbea587cb6a1df1bf0e9e2e75b8ba2d6117d4291edc58eb5aace1c4b9b6184028ba06ad774d47b0b6ce67c9ddbc0b22c19ed9e5e9370e5c62da8fce4e121ec13fd039236478ac9adb00f9ad81b499bff15a18bb191be4cfc27a68ef10908b3ac5f7119b436285bc3c9c88a03568c95ef6e5b1f3e3acf68bc297f4a8b81989ed48d9f9640c3ce3214e41b49a0756dc20dfb8833a8d9bba5dd06cd722cad3f99eb0e53fe1d52c70cb9ca7db0983a752c28f7cffa27a0c0495cb4f858a37ddf5a54a4a195322f5a8d2c84048c91cc67c1510f7aefc6010af501f5bef73ec02fe7da8619c991dac799eeb322117062d48c7e7c7cf987d12c838925dadd8f42e7abff01547dd952e40257583e368e72b5c138ebe37eec9d2e241c7950a8da8a8b216e85aec8caddd2af0708559012d6f5eac223007bf4edce2300bb4589a6149a62dad4204c13b81394b60350fddb07eac7e8699d0bdf4e10794289b3e466df9aed5de185325a83bdcb2b30a554bc7ef02f8b6e2f100b76b8eb3dec5016ac71c759a222e0cfba57fc6f3f14d1e987d2dd076cf6645cdf868417fb3d116a29234ae1559eb737287fb69ea8d5142969f595350ccb74acb847a4b0fd36cfb1f2b2bd77268d9add5fb2c48e799715215e866b11bdaa0f68c199c7c0eeca3d5db3ec80e66312868add323b9e54651a4fdaedbcfa157c8b12a24d6c88fcfb073113403b6346b2a5134ae87a64469cbe0f912ee1a86844defb769a33ad825104e26b2d56e296dd239ca66d26d5358f83a22f454af211a42e726d377ddefc21dbd8db4e91221faae31d49f1e285b7428ea45fbb11654202588a4fdbcbea793d6bb644cad87558ae015925da5c458c8838567f89c6f71cb24160c06b83b4b1a347a8532e94d9de3d39b20048c3cdcb9f98c66dc1a9f90c201459be662096537a10de87ebb299d19a510700bf1caf3f0d21b95b24448187b8867e0e92827dbdc5add21d3415ed10764f6ce086bb34806becca4463f4d94b6e08c108d339d8ce162bd90e20d4639f0a6431768ee063d9b1e0dff82834fcd021b58e0f6b507f50928dda54676c243b3ec8d91a4edc0a02c980b4a094d958a5b5ea294a93afcc3c8b8cea1dc1476e722d413fc4834e976bf8ec2e14351a8ff837d3de1789d7a7aa152264476df85b95bca54371515014b54adf632b85005c7d9845623ec9cd8dba5fdbece543b620be97ca16202e385d727d51d6765c04436c445f8937b7e8d630836cf1a816461adc9dfbb2cad27e0fbb9455a9aefeafad9f0c8b3361639a73cd799b9b623ebe57d1de4fbf714f4185d6477b53b6b6f624d84bf3227c059699fb942bf57af8f15f8fc8e72e5bc64674b9997bab9c1846261b9c59ed38931c6cf71b3c15b3aa4fd0194b1dbb09a05e19b851ce569394fe44b5c725c5e0d00f886f22c33ff2984074ac2c35223a19b9ebb3c06f0194259723a6acc76f05d5c27fc8a1d5cc559b8f83b16b002b1289433c316e2373d99b809aec928927cfeed79e4b7cf222463e6b77c77af782c6ed4ebd37ddc9df311c930e87a92f74f5c516609792d0d03ffa8b6ddc42df1bc654ecb2707aba1f3ad3d90108a4ac41540421ce65a9c00047c3f969002a7deb2b2b9ca8084f5f5f937c250b509dacbfddec088581d03019cc47e9b213d71589e78f4308e40a9caad9e607adfa3ab395d7d2cb94993b61470f3acfac955cb80e64890a5f7991fc7c4d73637c32f2e9f23009e1e7852ff2e671d31aea25678050b9f611dcacf9d6c3fcc6c3d94f5afc7ed38273af96c5fa2fbb9f0bea557c7000f84d2e792d20beff8d0206235c77b4c74071f8e8d6a972e8b1e914ba70059ebcb3883ea765263f3a746be7e59cebae341987bb5eb282dc4f6130da66a5fed586c6569281fc344ebae3aa278ab1c25ca8403aad378708d7a170410f397b3186d99ee770d4cdb3325aff5cee125cb273671ebdc10942f7d5acb38b9c5c209ca233f3a0c1392f4a2f508dfe86433b7486bc4eb29886db700e256aa0711ffd48b778137c57f4ae4b3328f6f3798adbd2fe87575faa51d07e8efefe9aa98e68ca2e2936dd5478d71d880617ff29e36abb4f331e65558e85f9537f891a5ae8be5324a7d12d70c1ff03ff366010e26a78bc0d3a202c42b5169abb9ba6b0926c42a7e709be64b24ad0156998e805111e44af5fd6c9dbb3ca1f8e7a724dc07ff0ca1d531c3005a0ffe6e0d0ec3468c14e03db1c005d8c0494efd4862410b54779c0e2c6a9a1c6ec9901daf4e6cbb2b0f41f93a24cea550b90ffdb9299317e7e2c135d9cff033f4c7a5f09035239bb9251fb77071a7b2dab97bb76de278ad4c4d0e10950b91fca6657fde7eb78ec3a28ebe8022a13699e3e627eeb4b261a1ad5a270fec02326df3132ed914279cf17889e5617a8f0b70af1bb5d4469052c5f4cf22171dbf158451c82bbbe3beaf307168cbcb80c921a9497d8d9f4c6a5e99fa2aed2f7a0c81b6b1c35a8ca0deff1f917d738a248f25512d5fee9aaa23e87aaf26b6f9be13578c9a935ff488dc47ae9199d14bde915f6d338b48ed87a109850c643730b1c990f7c121a39c0f219e218de7dd7307b23a22dddafe1891b71b3af641a43db492fa3c25479655d1a1cebb7d1db52ef3e5a7916f1074a4306b1d6fbec432f3c90b5bcfffe78712e677d44030e11764bd477cf187b8cc60555a14f546c595e776cc8940e00465144a7bbf3a95872517580be7bee8b9715d9f2b1e22725dfe0221101ddbbfd54350c729a04cfe0a7883ec01d216d63bccc68dae15981f7a5a2b1fcf2888aa3fde7eab1ae210fe2b7aa47b86571954e9152b5a6af0f19380bf5ab30b8b6638da0cab8d5735fcd3c3722e8e0c56082ee59eeaa30da1127b766cc9e44fdaba93ecf81dbb21c21542c93f966a5bfe7fe1e3bdae57302a873b5430af85d1848543dbab3b64bb9950177c4ab337ecee86183bcef3400f722ca56732b2db5470581882dd601c551163006d3e856cece345e5ad00dd4afe6ea7330473ae9f6bbcf11fda8c9dd93ecb5c527cb8d'},
	]
	c := new_context(.shake_128f)
	for item in tests {
		m := hex.decode(item.m)!
		skseed := hex.decode(item.skseed)!
		pkseed := hex.decode(item.pkseed)!
		pkroot := hex.decode(item.pkroot)!
		expect_sig := hex.decode(item.expect_sig)!

		// we dont support for 4-bytes of idxtreehigh, so we discard it
		// idxtree := u64(item.idxtreemid) << 32 | u32(item.idxtreelow)
		mut idxtree := TreeIndex{
			hi: item.idxtreehigh
			mi: item.idxtreemid
			lo: item.idxtreelow
		}
		// ht_sign(c &Context, m []u8, skseed []u8, pkseed []u8, idxtree_ TreeIndex, idxleaf_ u32) !&HypertreeSignature
		htsig := ht_sign(c, m, skseed, pkseed, mut idxtree, item.idxleaf)!
		assert htsig.bytes() == expect_sig

		// ht_verify(c &Context, m []u8, sight &HypertreeSignature, pkseed []u8, idxtree_ TreeIndex, idxleaf_ u32, pkroot []u8) !bool
		assert ht_verify(c, m, htsig, pkseed, mut idxtree, item.idxleaf, pkroot)!
	}
}
