// Copyright © 2024 blackshirt.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
//
// Test for SLH-DSA Signature generation
// The test materials was taken partially from FIPS 205 sigGen test vector
module pslhdsa

import encoding.hex

fn test_siggen_nondeterministic_external_pure() ! {
	// "tgid": 37,
	// "testtype": "AFT",
	// "parameterset": "SLH-DSA-SHA2-128f",
	// "deterministic": false,
	// "signatureinterface": "external",
	// "prehash": "pure",
	// "tests": [
	// {
	// "tcid": 313,
	// "deferred": false,
	// "sk": "198276F1CAF3AE81992E53BF1EC51AB370E74A22E27CAAE9B0C953B2CDF36B04EE9E93E95DC14F02AF76FBBF312BCC5AD207561EA17CB649E4CB3FA0AF5F5C10",
	// "pk": "EE9E93E95DC14F02AF76FBBF312BCC5AD207561EA17CB649E4CB3FA0AF5F5C10",
	// "additionalrandomness": "201FFEE926EBA71B8222D98CB8CC6BCB",
	// "message": "C09D602B21F3A0B10E4BAB37376E819F1E04783B8BDD4481FA9BE228B2B33F3686097B0B414C51CB51ACC480526CD8A23A91964B84567B3CA8A27873BEF15DD2CCFDA40F10BC31B54FFC920719ED23720FA11A10860B342B188BC77202A1C7E3B3DE6D75DFE74355A21C57B88194C870147A1586D511B0397283F65411D3D1A7B5149CE15D38EC2527EF223745A6AE0FE0D946D3497DF750BFCBADCC0C6B44C4539D5F30A4A8495B4E5E03CC617005204F03BF569825441545408AA6933B842ABC83A74AC7FE13A02FDEF98E923C904971410790960048FBE8272FB748783A47ED9509F2BA776157945556E0202D3C74F7D21FCD8271C0C57662C22955A8F685BF19BBCEB1881C900E8A0257C6BE5DAA50855F3FFEF961A964BA7AD70870E197AD1C9F7DD78DFA57121DC7E41A2580F039CA9A373FA3A25E97935CACDF2EAED66E1D7C46AE9674EBBC9FE2A158F93CC0665905B6474FB429634E144C78B7F6F4BE20DD57E6E74A3E80E187F4CD05ADACDFD463D5236CF64C74632DF9D5F5CD4493AFA705A51B95CA2F28233D9C288C9047E94145FB89A3652683737CB17A67A31F231C5A96F496201A5E5FC7D21CD0E7DFDE733D99EC67B0093DFA3C3CB0298FEFF55A6C106C6FBA26DA316239ADA220BFAF2CDA09579979902CC605AFBDFB4CC19974753D90970BB97C943265F7DDD042A9F938FCEB29646B97FCA7772837BB0D975A167DE5CAB9E728C632BC04118CD43D2EE67908E31CB0F25A08497E337FAF51377684B10D70907240E007D957C69F4625ABA8E60D450EDEC88B565A2B2808CD0C13CAB0D2FAE9D6CC864DF2FA787DB16274A73C4DBB64022757ABF6465DF88ED20252D47702BACDE7F5A27147353573829DB823B7DBD05EE842B38DC7D0CB6FF8952830EC004E1A985E171D1A4D45DAE572C712CCF024FA333ED5C61D532BFF12BCBE8D101BE64AAF8414DBD6039DBD08D0E1F3CFDD2BB723384BD24AFE9FAD3AED20B70A4DAAC66597F0F8A747337F101FC4BC0066ED3374C9DBBBE14CE19F7CBC230982ADDDCD8CE259BD11A080FEF32D1E2C9E1C695DF7A365E81B37A8BF540198284526AD2F4B62D86AC3E4D7D9B2F6F28A0B36A115E469302FDC2930654C1DA2E87932F4E6B829623F314EC627D342114B9DF5DCF6E9125B3A0D6558AEA20AB88A0CAB1CC342907FE82C8B273FA33D9535D7D26F04A7AE9396F6367737118FCA598D6A656878E91E0DF984A57DA85171849C6A3D6D6346F5721494AD609D796CD208D09115C231A0143FD34A9D21A72AA39715B07E61D3291F7F289A18FE5EE04421C725D2F508994DE99E408D65759BAEADABBE7EBD8E992EA3871D5C7E89B38061B012BC56D74F55936D0CFB01CDA79D8419A2B1DE41F434837BAA445E2DBAF599425A0D121FC74F5C9CC0B1C31DA94DCC7B89397F4DC2BCBD25DC1D27ABF2541FCF18AB1B73180E5222FEA1FDB25A6099D1F05081DAC5B2ED76802B2D1A725B3EBE641D7D431FBCCC0B1345FFB0323E510A389907301384ED95EE3A30E5196668FE5130F1AC6AD16BF881955EB348DBB0B0114780DA598FEE56C9E7148AB54DA072F8478BE2EF6251B87461C001DAB77D02C4E533B9D96045DD12E10EBB8ADF594196396AC5DE75964400593B9F6C0137D8A39E690E8F37AC630D6A5885A65212AF002C03118F21A12EF4C2F185C452476A66B50D9C8E5A6E994AFAE77FA48A07F2DEFFF2B46C9E8DB13BF869FDD1F65DF4EAFC10AE44F1AFF2E06FAF1DD2DC275DC0C27C224731677763518D3E4C4F09FA17B95CCCE7C7B45A2239E5D315F102C937B54DDAF175AE47C8F776F84CD12CC642C50FD5A65F130D9C6D97F578306FD94ADA0F79154BBF278E022BFAD551C8BA2F5E0384CB4DA3472F6226B19C3D49F4F24B4A148B5B254649DA2349A64270C31E3432C224612594EE9BD43B920901B14CD13C4614E6EE612127E6F1E292E2039DB8BA9EEF96C52F915EFB7ABC466E30CB05DB89450E7BD8D32158EA91B7F3EA1591810039CDB7285A82548FBFC1837A1177A8D67CF8941FB8F36CA6BE20B1E5EEBB3C40C17FA874DC5881D92D34CC3FC8170A429DE1A552D14380E1419380DC5B82C38C014B911CBA45B7224B656238D5AE3A3EFC0D68B2483D8C529C62B9937ACC3F906CA2EE035607500594EE905D961C44FB27FBA99B12302FEF4FE7230B4A4C10DBC2F8551AA96239A5A87AE3772DDB3ABF6D04E08BA80289C1BC976590ACF87F7765BD38D0DBB2FF0786519D9BF2EC87B477D004CAC37699FBC930CCA86AC0F74516D563B490B28F71CEA30141FD52F28940D050A43E954CC972C8836B24CDAB87929BEEE575C885C87442600F400BC44D9CF176154889E104BAD97D157B04B42EB3414CC2A08F7AB7E5982D1F9A07A3EFDEFF70D9FC5EC9DF5D8E74F07F6A60A162FB17E3FBA34C0CCA737311683F932FCAFC80DCA61729CA244865EC9C452A59A9955F2E366DEC5EDB16F02628EE27C37B1035A9C40A37C1294E51E7012723BB999CFF8F020E40FFA644E7DDD9521976306714BF00C3F6A925623C776D92A3C2F4CA794264572B8FD0366DBAB45D2466C5BE7AA5EA178612DE63E72E9E103613FF9B3BFDB9DE34AA0DFED786D5D50C0D90DB88A4A6A35D2FC832209802388EA8BD4390C06AB4414D62204847474E44FFFCEA672DB9F3568F5BA5B2FA2C97CB55461FD51AD408F7F7084197FD33B9D57A2C4C30CE8ED4C7925D64C961AC4A8EFA1D7B011DC9714C2CB8F5018086B4F425075E45BB92E9D1473C9E8B2035AFED0AC21DB128DEDDD97108C2B7601C0330E885FF119A545018CFA4DFFAA2E354EF70551E84B69C7A2419F9990CAAB8762736416E75251F432846D44EA303F6D20B146D70D6433A7157FB2431DD7D97ED1D47E3F075EE685CE02C61BE28F476494AD617A398D6BD0A26B65DDD82006F8A05FD42194D40A922B70546934E6028B4D8A6324D079CEA5F6030301F11206227C0B01E51A84EF07C241F4082361D3B57D66FFDE4282F3A234EEB673DBDCE41F8887CB189B7FE23D68B5A7D42C0394AC86EEEED5318EAA47139D64FCC257BD7A26100BC81E6A945C3C216CFCDA173FA9EB78DB99470A3F844FD9832FDC2E6EC5A271FB6BBD7025527835DF6102FA2096CD411B212D6FEC117BB93833CD0C821B927FE6FABE0CEB06A9F8F9331BAB4D881D403C6E39F145997CA9689886DF5B7168FB1C50824DE6F9AF5522630968CAD451CF13287DFB06AEC0693895069A5BDC6C029BE68F9F473068BA5930900602B54E6F22D2ABC77404D19BEFC97E5FB40885C2791C1E19438491CEEFF20FD83AB032B6E4BA92E19ED51EB9FFD313E8FF58AC6918DAB6456C3329C5B44AAC82BEC16F03A26DA85061AE9D2F517A5C7D4A56098C74CEA9A9B3E5149D0AF4803C0460344C405E3EF8E52127B2746A2A80D034BA4486A0F2E31DAF51E1669D71896111997C0B2CA1F4AA803D77B1B75915D67B2A8C8DF15D9DEC3F68F252E9891298D979CD8FF10BFAB14845D44EDF227691B4DAEFB00A62DAEF197D0717634CE0647C46D43DFACAA16ADA96E0DC4CB7693680559FD9ED9EDFADA7C84AA266D548291210F6485906F744A4CD4EEA0082A7641F6DFCBB760275728F3D34E21F46382970F16EE41B88A47D0105DC63116EDAECAA69E89EFEC92A710511C10D83F85A71306058EB7F51CE080CEB7490838A94503AC8EA79B76889D9ECDE45E980A16885A65FFDA5CF15B584D3A0078893075F4AFB51AEFC8DF0D12E16280124E691A804641797D2D59FA1E9B5686A98969FF1EE032C7B38B5DC9D3E32C335610F6AFD3E389E1894E55277768A64C91B3F03E14B99009FD3DFE0928CAC8D354D063C4E7E83A99C77EB8AFE93004B19585949CB68003BAD4DE970E7C516041FD3F577B193BD2264FA7BF187365E7954B7B5B880CC613AC4B7DFFB90E8A4087972B14D1C54F2CF00EA063C92D4F37D498A698BDD8F76C12101DCB462BE0C6B271EC68AA3A7F3CE338348079D923C917C32B9AD53DB17400D54E50013365248F193CEDF667FA00327CD56F4DF84261611FFEAB4F6FE0EF5EE3D0A43AB1B8B8A88179BB3A85E8166F7B0AB62C1057D07A8902BAEC0DA508D57673DF7D697B3C320180A5C8BDEA64D9EBB9F578B665D2C24E0EB5EEEBBA2826427824EAC2012870826C91E31A1E893EF1A5A636CC4A4E9A5EA27F92EBBF9F9363BFE74629567F91EFC2C304003064CDA1A1AD8A4D8CE629BF4D4041931832457191147FEC2BE09F30F3C3B3740EE89EE313AB1E051124783FD47109F5B085B3753713E8CF48E04CBFB39C720426FE315635F219CBA87D847AE3C8CD779F52CC66C8D9733F3FD4D62C77C682969F5B08A2E9A9477CEB7B4EAA5228A31E0CC486353211602EA01AFF7D6E0447F728D7A286E7DA3C2688FF772807135A3F514430BEBDAB6D41E1EF7C25CFD07B63A456BEAC67F5633D8243E19F53421D1D40CF4DEA68EB4DE6840A7B4B18BE6A699ECB6A25309A0E9F2F99AA0B91F14B5D3A95E439391A2E0F7CEE47769493D72D4F72919FA058B22508860597FACAD5CC8010DEEFECB9DC2F6A0A7DE2BF17263530A5D567BDCC6E1985D0F2154A991AF9D1078DBAC808D224D94E6B0E7137F5FB9C4F3014C4A6D30DCBA7F8BEDEB57ED519EF19B512C28561BA990D91D939C07D8FD1CBC86E33E9EBBDA07D4D698CBEE7E0454832B485CC67189F48AD9291AE49F5624B9C9D5E1A6121CE3BDF2A9D000246A0238882B6DFDB6D682789940AB9F880A8EB6A8F058703CDCAE894603AD04028DDB84C8A2EF1E1CCDAA12562E72C0A629B1AFADE29DFFEECADB67497ACB50F8E8A71C1151C949AA2CA936E0374B0833F804016495ECA9A9ECD681EC994AB6049A599136B6B8AA3B26459A9C37ECB55CC7F08420CFFB4279DDD2D9FC046FFFC7356EDCFC97D0347C24D15FE866877CB6C2965C8901FB7367563906FB34DF1C763DF123A4A387E32489961C4352A8B2E4CE0ECB10E62DB8591370847AF4BE024124B291196C4AC59DA742A6BA4486D7DAB3FBB947103128CF0A8FEF69158A67204060CA3A8366E08755EB421EFCB2E902D99A055BEE52B1FEED14704CC21B78F951937D3D89B174C957A7A9D22005E37ADCB1849E83B8C3CD9E53EBF820382EFFBD7214D03DC5B46E389914B2104042C90C9084F11B366B7663AAF34E1FBD526C59CA1272DEF01B61A29FD4FF3F37688191FBA572A488B9DFE4F3C0492756FE1D8843F988D1E4C4B2133979D516506A33F41A951DCADAB05352F45793A23E9B1C74FB4F996B6C9C3709705D64DC1CD44C877287B2737308C7ED64F57E1BCE32709E45E1EA9CF1A67BDD0880C3A29DB848627361E4AF296256D5DC8B01D8793F9A340FF2845536BFE95726EBD5C9EEA46876CDE75B68768080DA37215CDAFDA2B8DE4AA257062F1659DECA5B2FBA3C9E0739660F7B221DE4E656F8A36B808EB3A256A60267E5DDDE764919794D6CE7897DA2B1EB9E9FF96EE0B29834D4956F634807B80743BA30B914F4AF74910E978E9BDD48CAF3D6CB5A6DF9CC98AEE2D315CDAA77D4EB7356C67DA5B259FA6758AD4B3727A7AB2D1DBFEC938AAA70AE6EC75E99EBE9BBE2C5B374F3F80196B7FDE8943D471DBA21AFB99423B7A126DBBA65B74901E85FECEA9254E1C95AD6A1E3A444A1762B14261050823BD696751A954E5EDEB37A5C329A1A685B33DA7231E57ACA3CBBBC2A09347AC36E2AEA0742FD88BC4B8CCC2CADE0F06D90245890E3BEAD25DDE972A35199DBAAD0283D3307BA9CB3D4CE30DF1B58A3AF6F0DB3E4EF5AFB9B5DF1B1DFA15D8A8C6BE77551806F7B541937EBEF59FB178FB91400DC1647825579CD92730EA5EBB0AD9ACA32E86CC36FD9CA2C71A07568E074B0759D1E2817262A5DBE43CF551E35A99C54C2EB8C403EA11EF42D7DBCA3381151D82CDB955D025DB5CF289B648EDDE79A2E53AD7A424CDD51226B3A64EBE98659B84E3305CFD7E0024D3DD92D8FC38A3E9259A63981C9A00B329B6D3D149AE3A8462B38090C89E3C48D3F43F2580FFC8FA84F0FDF91CC84F0574F8FA39C7D318120213D8C53327D922937F606B9F75AB24EF9BA562C03D973A78B4B8A1C0CFC83360DE9A2C23B8952952BD36B403C7B92C9ABB098F0779F09D3FFB7DC9512BE0C934633358A145E0F92AACDBB1DAD736F67D0ACCA198FD9794373C7204B1C0D62E6F108C3ABE3637675DA28C9E0D28D9B2002E8A285950D9C19DF28FD9AC3D9BB74BE9DAB48A3725073226F172BE3486C6151F424C7821174AC41671E33D6A8D4E144BD394EEEFD2437B0249719A9ED80FD6CC433A8CB0031E7DC9A45C7AA10A7C978C1196435C93595ACFFC7C4094136873EC8447E625DB25E216F082482C12787E8A06AD074BFB5B142A6068D5E5356E4BEC888D1988069D3A18E23EB7A783BA37D26175035E55FC799ED0EDC3153EC455A829CCE74A4AE0FF090C5D4774F9E417237D14A98B1675B970D7646906A7467629B3B18C9BDEB4E70B001AD30F6C500239F46A5BB4ED0859B667C5FE32EB0023E06CB4C4FC1E0C8ED9C99793702B2136D6965407CA27E2DD77ADABA76D8DB1A2948AFF30A226998EFB348397CB8007620F328CE38D94AEE09C56EB95AD07C35C616314788D3069627AE29C78077F34624359AF30EA1205A8038D600B89137197AD8A1700E24ABBBE6376F5933DB16EFD6274A91F9F70E77863F7C248EECCD96F76D929757C96D6EC784EA0D18A699FC6D64ED76283E871D6009497B937330D044880FDDD77444C3AD72C071147E70CFBB0F97CFBD022F074B6A0BAC8D1AE187F60E8B9976550C0524AA885735C2877BB5D68674FB26DEC0118632D379796E25CA06339BEA3696418492E69BD2309D7E4D8525FB40AB9E39AA65C01C9690A81B365A87C340C4F0DBC1C72099507935E1A2C9641184A48051D98460EB026818A53C471508223047B196BA9FC0FD67BE1B50D284AF45D4524B52BA038886978661981DF11E9486B42778B9E5E6EFE30BDD0CF78298C9A0C33D55A98ED657C06B8CA18FB3F944CB02D37B4E500901B7F4E1805B48E22427E15C1735D9976A3F75D8B2F7AEE4D49C3855D9B6C0BB0CDA633F30E915CD991E74406488857D10EC8A4C095CE374E725DAA628E200A87855D4ACB2FA73F47B7F35A66C961AAF325147EA5F4900D1872629B4DD814CCEC4E0D67F27C7DE58C6E9850A3E6A9B10EAA83765B0C5895ED50C6481434ADE00796400F7A6F54769C6F8AFE897D5EDEBA77D0FBB91C632C5D87D747F21954176C21CE01C46328DFA53C92BE39B61DC498B962694C1A02D6980573A24EFAB22F2DC4B4A642F6971CE11C15BBF2FC32D12A2642A54882DB21C810F85C8009FBBBF784BA6B8747EBDA5EABEC273BCAE69161F4AC4AB6AAB4E8303CEE2DD1F5C7CD445086D98D94C5D670F84FFD6B0B5DB63DC95248D73F0B7D5E47004D1E5BD3ADA857339981245AB33C8389C2271230308A0C88A4A36F2578E907FEE748025AFABA770F9B3CE8C2C66DF5B8FDB7F5845C2F485078558E24B7F3708143EBC8A9F48040B7AC6E5F78DA84DE32C72719E86A4AE9AFF1F7DA3A72237EFBB4C247A5A0BDDF169F60CF45DE39475390004835EE24448B906866D497E0177CB43EB221D86E32105D070CAED67A1758CB721B8A9F323967E41F13D2CD3C1EAC0FA5C0F69112C5AB8AE768288B28AAA43A3311B58C2721743544349D1ABCF8C53098D7801F528CDC27A8B1C1A76FAB19BC2E8FC5024E45E726DF491DEFEC543BA90F97374267D3CAF91303D20E48537F62248A6EF8A1D5C7D019E7F21D85F02B7ABF09FBEE0D3D469D8867D81615010ED167A3E018CEFBB30B86457FAE705260EC1AE70F5625E60504A23DF354E04E1599966370E6DC4562CE5F21D41342E9DA7CBBB8642B9AA435D789BC5D30CA132C5B59C2974BCE1CA47F13AAFA5ABD8FC1006EBE670CA96E5C2DAF3E0281C475795A7B92A303E9483A23C50E9AF7D1E4168C3E22A5436DA7EDFCC581940940698DADA1CC3FD31CFF221301D5B4976B21AE434842EB52221A26BB66BF020C5C3BF879A5051880285ECF2974C85D946354BCC88DF14538E333B2B94C6732EB2897DB5F6917EB27E93C358D7BCE85D4D4732398AB2BA4389B6291912D02BD5DEB4BF8FA9C310786EC68F3312AE09B75C4DFBB0AC51D3720927891719ED88FDC6E5F6D17434AB48F7DE8B6E34B36B12CD32F69BCDE2BBD59623C4451C1856FA24B3F68DB0D6EA52E9C9A3583779A5CD7CA53F60D7ADB1CD63B7A85E878502AB36C2D7DA80D7C7FC93DE497FB02F9D4E825BDA2EC38DBD0C8E775588C38E2123495377C4C8281946C3F2FE84BA3044C9307BECB8B85C0EBE879FF2AA2E9BFF9252F3BFF4E8DDCA6F04827AC24C44AC81217414C3108426F94860A282972DD94EC53AC956C1663D554EFD3CDF55471F3A2299C7F7DAB4CD2C5A715B2623096C3161C0195B7ECF1AE97BFF87DDA0717AA386C59BF35F3B1EDE864825DC5FB944C6DAED40CFFA960FBE8D1732F9934374805DAADF77D0471EA29003F17E8DA800AEE92B2114F1D85E564D7C4A7DEDBEE277B6B38460583DF20BF242A848FC4D3AD79510A885CB2B33E21B37A5D24310F5385CEDBBB87F95CF91A0FC4035BA699DE34E9D8ED2F73F65727C040627CFA308427852A29A30796513F39FC530ADAFE6115F75755B536D9B0F87EC31D4B9B331762CEDD5908AFD58B3E8E240823EED6EADD8BFDAF11925205DE32D87892D4DF63412042E0C5DBED13A668E7083CB7E3D0F756F22AFE7537A4AEA335F5C27CF4259660BF07BFCD40D0B6FC24493701A813279AF587FA76C4012701AD05ABA30FCBB21F0AE4CB0B6BEDDDECA1C3765FA65CA8E198D148A645A1458B122ABB1EBC57BF9BA8DD5E51F5C06C3E2E3F17098D392B692368FACF675AFD6936C0CBD72B0B2CB8CC0498D1C6CC4993A0AF01420A7B4CDD02E629E80F8CA041AF241E3E530DED2F822184DA172D504D500A5B079BAC8D54FF1FE5193BAEDA51DEB0FF161A9A9DFCB69DEF97D04CFCE7006596EADD7EF1AE3A39D9F109A4CC71B95426141450B3E7F438858D5BC88DD810EEBD081F93A604C41466CD8292343C2A4A605D250DD5BD6DB67D8383B5C3A0065B833EE1F7BB19B24B21EA0D209E72BC09431E699434942D9EFFDBAD5950E5FF74EE2005F1466D68C9F259A1035C6D922BDCD49BC215F57C892F276524E2A5A4C2EE6A8D319D99DDDEE07E8AB01D5CC5650090FEF5A8EDDE7C51A28A234C49477C09BE6022D292BBDBC943AFF371CE2BB94AB16D2A22AE814E8D60C35874A6219071FB7E491610176DBA20A3293B6BDC15FBFECA6ED9B97888077733E90075FC6C6DEB5F4EE326B8152046E39B3689C5C04AC4CE70138F7BD14A626FCF2637B49EBCDAB3002C27D9C96EDEFD548AC3EA77465921B514B84721EB8B75BDF027F31E9B6E5E20010B1A6B79E2285AB0675DBF1F60F61955500C1AFBB50C469252AC9739AEBBE78209D83C73760521D242D6F8D208109CBF2CCC5656E12ADA488DE17E03FB9D865F2FC72FFDB54621A663FB258F54D474D1AF93D6351A174A39D5F2BA98AC84CD68654DA67CE14C520301716D2B64B03A477A2A88C905ECACD544114907492318D1278A3F8F1CEEFC375CDB21C7EC8F4A1FF904BBC455F4F2A5DCC26ADD84AEDE22395ABAAFCF344C35EFDDBDF7918998AFEECEB52846522BE1390FC36823EB151AD2B250843E39EDAF2C011681D62BB4A02A8EC999C8B1D58ADFF9E9BDE47836065E94224529C23EB8677ED91BDC0ADB22CCA7E05AF174AEF5F879477CF1552D061DF28CB14E81470BE9BA0D77A7CE032675DB13117F54F9EA4671C671CE277375F580EAE03150FDE0B960AEEB5FF466BFEB15A464CB238707D2BE024B61016B98A66D6B0D8DEF3C193FDF35065BCCA948BC28723AC019E3618E77CF6E6A3DBFEE670AB7083D23E85D50647EAE84167FA22C6C8921F0D3A25D75A931754C8D7EBD8DB91DDA6ED5B54549630D6376580AC0ED1BFBE8FB4DA884E425DEF26832C05DC8F4078ED66CBD2855846E98578782539C9AA80DEA46B29448F3472CFE0ACAB8FC64EAF9ACA65A9529E62FADE1F0782B51DCFD33EABDC2B3EDB3353102E70F84325089CFB3D43099CD92CAACF9A0487E244A140E8FFC0885349ECEDC402728F493294E2A6F9C7665EA8C2FF343F651BC8F75582BDCA3AE807AF86C293A1B26FD850EA34B5CD7F37D75F0B13D7D837EA0C709F76625AE023674AA01621AEB569CCAAD76C29619C587DB7DD9DFD9222B7C5B871491B7F0AAFCD03964215FCFFB4ECF8B5FA8FFDA27DC9AAF56CFAAD270D8CB6132163926272A55769CBEF55F37324D84B24AFBF6DD8E9D4EB7DE1AFF726CF85A80960249D281D55B9FDD69C52B518E70CF1D3F69334CF8345F0CA8FC85F453068320B0C5A31CA1F1B32E43D6C3FC5B5FDB9FF4C6737C7B315CA5657473898AE2B32DC186B06910C3E4B3E5AE7E54DAC4811B860FD7073345A7612FB4DF86A599DCC12A9EC1DC7B61AFCBCEA6C122938B5944FB182266A4DECB83622CCBC08EB359A6D011E034097C34A8767BE6FEC9098DFA746D39FE40ADD20BD2CB59B00A2646B5A48B2B2086CEB23517621476E99D4FBBDCD6E6D468FE31FC326603BCB24C0B8AF2D09C18C56AD15B42A2FD72A90471D5880BFC16B1388541A3F18B582AF5D714D4BD7B5B73D7C7D9EC970CED3FD5EDBDBE2DB18960E0486D2B0FF08C43BEF34F8F3C4797C2300339945DF6F9A6B0",
	// "context": "DE4E64C30CF4AA6C889FCD8B8C29D5C4DA1607B720FBFA7BDE4E1C5D5B733CAA55F4AF139B88C627D61EE5206786699E7F3400F576C0BF8E62004CD21C818A6EC03411F6C855F8DA0B7E78DF8A5C7B2A2038DEE5E2FDDF67EA78689463D1A54FFE6F7DE3B08AD75E1AE2F25528AA07CA94AFA4C2D089DD3E18C280A0B313BDFDD4A08A912710DAC4FAAE6FBF3BF72A6B191CA721CE7AEF8801A4F38B4FD20D89A22E4D521520E73BD0723CBF12DFE30C4ECF72",
	// "hashalg": "none",
	// "signature": "45F33C1F0DF0CFA587FEBE231394E160199EE47CA8819C82E21CCDEC53809A0DC3320B66D8F29FC294D87D0389AA6E25B375D245B20B16816F0739CD9FFE863A259CB9331AB93E3BFE70636955F352EDEA292B8CF25A8B865747B81FEA73B2F9C24937CBED62E479D654C3F1817F6EDBAE2B67EF845681A645A55B943F9A566616174E4698415127D5C8CB88D6D7311132E62D0F335B1F7226B787B0E4E45A9C2E4D93AB0C93F18FB0F0695DADF897D76187AEB2ED55A28A43BA7ED58CB0D64A09DCB70DDCAAD472B69B57949242A8569E4C732C716D07D341D634BEE84CFCF93C3EB100FF1CB6FF1F64BE283AAF4C4B842F0EFB24CA24DC244A70A7D8D9F231648B6BCA0E2E747A40E10F57D838048694033F24761FEB635BAE07C5E954D67D1EA5A243DDE59E1028E7FE125D1C29BA4F472F0788EA871CFEC58B854E487E8178BE8E0A22056E346F3CAF30BFAD0429E4E8B115ABAB3D7B8653BE2D12D0F7F41B2B2633410E3E995C3BA5437E4B883DC7B85FF4B1ADE28460FAB4D471FFF6B5EBE58670F405EA69B4D962D358C05950F67C70D661142020426DC32024E0A7CD379D08295944A5A7BE1B97C72A4849CBB916E2CF3B180E302F13EBACC829989DB86418B0D8BB2C897DB2006ED4B5D69C6DAC5E603937897F53D62666BDF30EF9231D6BFCBFD4C5AF57C77A7656D8B2E15A7B13E8277B8BE6DC16D744A465CB81A10CC766A8BE2CEFE5532213B3EA6EFD884214637ECABEB9F966699A69163A51F5661C6B830A0ADD66E3B931787D0366A4D473DBE69A4063C1B4EE8BC9E13CA1621ECD4EA78CA2168C96710BFD67D7D972714780899B71DD35AB693377C2521E73D6995A884E606E94407EA2B4B2ACD16C8C5FA7755224225E3C25CED4065FE5B1B5C343057A3793300C92F9A8F93F3E326C2E9BDE569E26749D5E601ADB3AAB673C3B5F54AE5AC0A8E67F30D0BC2EC144A20C45193D98F8F074FBF57986DDF71A1CA90166E9C3E07B64D280954CBEA0359BBA470DD7746F96B90990E51A47478EEB60210A44BEBA27C4AB27378143E029A55D8E83D24517D6882ED36ED833B85142B2F299CD1F8ACA9F0E144245FF409E9C09B32D1E6EECFDDF13F14FAC9E1D537C1C4B1063FEB0354DDA9D217687949EB933BF055D12BDFF4C9B9C162B805ECA8D63C868DB892248C4D1D844BC38939937CAECFE429904117D349F7414D24F7646D42FD47BE945F7EC6A3E6600C44D4339CA12DAF4D8B58A5437D90790C251A9DED082E7A39B305818991147598193C315D907CD7778D9EAA75875C2DA7F61ED5D1C2D5379A1BA7F23CA0165B2B3AD0C3D13FCF9C3B36C4863002FDF85884C3ECDC4BD9D39401162964C04ADA1B428B45866E2764655BF194E21C24607F120B56238A5479EE05DEB501BA09E714677C395AA5D1319D563EF981A753545ADA177E4B1A0F6A3B910E00EA6DBC636531EE88E068C229AB2AFDAD76DF51CF197DE702E081C786F18D9F28EEAD02B10D9DDF10967F8E64DEA3F51C4E72970E4FE28C361D893265FA22E573A4FE52154684191572E36000A758CFF2C459E23C9B9B1CA962DF4305E7C0789A2F00CF43A0F9E80A65D63B554F673BE96C6A36D671949BEA147A98AF4191BD8F61B4754039E8C7A3B3BDBF494368A556E49E1F0B4194E916B9D937579CC24C1ECD69FCA2ACCB0A8E63F13B1D6E1285402F72753672FC6A149D9FAE28FB7E90DBCEABD56993158F9ABDC2AD178D81296872CF444FAB021B1DBCDFC71AF3CE118ED7B4A8855D34E5EC5316C7EE7311327A28CBAF0B7190DA8C3C72DEB40D3DDF851D3E9240719074586A6FC0796882AD1EB5D1D7CCB3647F016CA91D7AEE1B6ACCC806D13F59A93D42CAB180682E4222E265CE90C09163CA03D6C63B2FBE8C53F542A6D8897E3D5C5B2EE781308668149CFAB81601498923B3356A1FC5E87ACD59205B3A789C488BEEBA5C4F2D1B70C8FC21154D4B6DC42CE16A93650F60F19D8D01593651BD60DAD6A1A3668E571344C3268F367A92521F383DE5F4A292A62C5031521FEE3E77C193CD8EFE5A4E69D5B7136E5E64A5C6EA6F53C3B3FEF95173282A673E54BAB8156CF459A6F92F75A3E14D62FCE2241172E25080E0225A6880967857BC058662EF1C7F9215080133151DCF7A897436606D53B2CD4904DA36A9146E833CD8F57847A7758498A6684EB4A99EAFC324B973268DD989E6DD73923A57D45A93FF16E2B7D92CA4EE484CAEC282A4B5CD59E0D559274327446376780BA0B4AD20024C0F1DB258A510D560294ED3A8504BDDAAC76A1BE72838BFC7D5779EB15D9A7D4E5CCF0057BB2124DB19EB737E7DD21F960B72CB3DC3FD90309C595A08E67D7B6207F067CD9D1EC23DF9B8EEE9DF2BA4E390DF6AC227926A73B78BFE02FCCE1E608AFE5DA2AF05C3A5BDD16966112724DFC32F6D32F6D39A026C8CEB56E347DAC45A3B1C0BECC0282F292A0B5ED2D36C706133D18AE2D252F8D9277C443134C78FF048167A3D1D94E0AA6C06B73EC7466CCC03528C9869B86A04EC51369EAA006BAE658FF49F597C72463EA8A8BEBE2BCD58C4D22951431B43C653C1EFFAEB01027FBC03A79FE7829F6B3B66A698D7396021BD92332EEA3D2DC485B1720B5BDB24341E75A676CD21BC650DC4D405D2557E874182BFE002A7EAC723565AA0FF2825019E93CDA672E13F26C6B1271C6A0F318BE29A9E1C2AD9893D2CECF135819D21C9A1C6A6C6568FB2C81EF15811DAB00718E8EB5C3C81C3E7842AA385068D12BFA5A952C84D00CC070DB07FFF3E5A9AEA57DA2D2FEDB95C1853216D4A17AC1F0C9D233B0B98397DE6264E90C96238EAB78FBEFA9699533B3B8B5AEDD59F1E603C3EE40F27FCAE578E982383D68C6936695B090A1545B1515D2DA5D66CA6FD80DDDBB73AB47C08771DF16E374755EAB703435CF049F4429BF7CC57698E5D674EB6423342B391C09903D4D82DCF52EF2CF339B5EBD8E948C69FB0E1CC71EED20E0F6F6A19E002F2DD727D0156FC3FFAAF9A8BD8D5BCC359A2144AEF4D7E78605891A7987FCDD59560F55E820E48405528D01215EC920273EDDEA684B01E383AD82FA3E139B3B946F5BC4AAEDBEE9755754D8C1909C4875F40EB846D9661D3857DE1DDBEE8DA72634915C286BC99654992511C8D756112D13001116E48ACAA952520415122D4D0232036AE605C73A262671E4AEE01B768E1B94D183BC5B06B64D3BF4B885CDFD13AA2299A853704F1C347F52B5ECAC30D97E6B0F4164EE9F4138F50BB03B31BE5E3535846AA4951B534265299A6CEA25C6F6017B1E50DA8360DBD347AFA0ABB2134E29C712750B74E7B232E8D7161658A78BFE2CA8CF08F55A90F90F8761DDEBE3CC78D07280F275BE9371678D5811798BDD7BF125C30675FEB868D7955B0229779EB83165FE5672A8F38100757105B337B7B2CD3D1D3201E71D0574D0EE8B219F92D1916BE2A4DC4347D0FD743B11153A00391E4411EB2B79FB5880F3B31A91B48C41FE1EF2C6F9D7B4D3B4E61C416C3656C50F422246AEF0253B917A34CF867FAD7D2FC8202D06EA7526B586B4E5B604A32F5B97170DA6A65103FA637A1B39F857414F7FDF9AF0CBF92FCB38DAEC89BE5D11328B9BD03E74827ED64289A56569A8F699DEB42D414A9F8DFA0CDC683D0A472F7CA0E84DD3D0E2473285EEBF55F696E7C26F88163CED91F5B2788563C04272DDF8F2409756461F4775E45FBEBC21AE145D22BACF71D630F53D41136FFB7DA0A55969859D3B76F87A214B2225A8DEBA0A9EABAB0C3FE895097A65F64F7661FD287CC52737D1A70E2D12150F2B79F42E9AC18B72F80BD0FBC5243F508F141F41A197FEEF24DF2644A82D66BBF4AB022756C33BD4F447081BC5D1416C138303E9D4D87AFF35E65CD76ACCD818229F99D169E2DB09FC9610066705CA25425BF7D3CA370709854B99E11B024F11A6560A3E0DD1E35E46EBA0A6F192F1D73F90697BCF8D9DC9735FF6FD5D492896121616653993ADD03CBA8E64FCA62CA61753E24FF35D210562E625DEBEAF7AA940E517FAA0CD51EBD9EEFC5DCF7F22B97F20F9570EBD34F35F3DB18A94DC11CB918F1B3B4BDDFBB78F50237427D7ED7309B2724D234E7EB632497C7C1939C05C0608087BC858744B0A1A837D62D057B6BAEE485C897143040BB5308D9077BDE0E8877A9B9B9892985FAA4A457DB8A320F42631516DCF746D3666683562629B76AB46500DC86E95785DFEA29962E6D21B39FA5E206C841575D8C79784C87519700C99D13812FAB43871CB0BD1A65242D0166D6313D87CCF8F268BCEB02D22CFFB683CE496499439C2DAA0705F612F0A7D61A8A04B41E528BC73E8A68F013B81E3E497327B7AA96D281D369D14758788D7A2B57567F3B95595C2960EE4597EC62F5F6F82DE7ACB34AFE2749AA6CFD4C26510F9DAA4750D4D95B37DA550AFA02D7D7ED8B522FE86C7212DCD55B7C45BC2387D4CA12F377FF01FBA6A5946A86FD192A7D88431409E6186F989E83C3429D1398586AF64826624988D48EB5D0F0990B5E0D1402C124C3CC5A84242B0FC487A13D197D8C5C560368B9729266CFF09C641FC9561B3F717DEDC8521F93936E08AD99203258E41DC9AB3C2339FBC919E0E0471AAD08DCB29FF6CAC5DE519D662307D21151D8796A3B0572D2BC9DAA8D565FE5B30649B2F66E5C6E18BBC7A0F48D507B5E93DDD9850BB6EF559CCDD40F7A8937166F75064253DA39E36916115B5618645E18C3973C5A5CD392963E393C803BE5845A06820EB8F8A1F9453BFFF7460F694EEEC9578E1808CC3BB7EB08E1F29D8261FEE147F5F7C94B65FDFE5F7FE2FEFB430BDF3A2417EEC2C406EAEAC70016FB860E505F5E44F67A3B5E14A395317AA256A84FC7609F570F3ACEFED41C934BF459B6FE5DDB39B5032FCE3715BA57C36CBB1968BB6C77C5369834BD9C3D5A9560595441E78831CC141AB7D80E290295230F1F4153B61E86430AEFE42EF6EABAB62188FB980269B72FD65929B5C4B893D11FB0F5F3D7CBEA475769DAB7AA9FA354B4E39C1FFEEA3A30E65A7B6997201266E90ECB5DC6819EDA816ADCA84EC739F0C188795E8A307636F848AAA715135C62D4CFC881358D34160E981F4EA7EF8C5A6D6254301863E86019EB4AC500259B5AD2DB169F322747DA3DA476FFC7C4E564E20710C111198A00ADA8D66C6947337C91F586402C73B9F1A147A98505CCF24823B9F7BA3BB55887682FB398616EBDF74C1D1A240D72624C43FE6A8E769D570AE5194CC59E60E3DB2416236187DD317F2DFC668EF4F23F9BE3831FED7B7A76345FDFB453B3631E236203A866508063C939FCACE9BC303F30A4C9BA76C12EB87921597CF53492686C233DC9EF45E293952A0836E1DAE197289F401AA581EC1AB52561A4F877B0BE1129BF1C9D088D4B1914C16276A6D9E618AD7414365A2719D0719F1EF8CCA60591DD23B18D9868F69324C485BDCC7393C2CDF2C634E29ED0A7192F7133990028333B7FCA8291EC220704027FBA21195F1FBC9640F4198B533A9793FAE53377B5307D6ED24EBAFBBC794059666692B08913018FA89422D6945FCF68383F4D2891E4085EBEFC8DE5B24A98664FA4425A1B62F2CCFF50CDFE81EEA6EA47636A41B82B292BC13997199FC088832545A23F7115737DCC903A07FC2BE52469C3C9512B46E42FEA096D4A485383E991860726A5AA11E91B8CC736D26378C74EE190C5186D030111332633DD4B9C630054B1289E887A683C45B775DB532A3B1C58741B80F4CAA232115B5BFE530DDA19C2FE84C19D5E31D7FF25D5F0A4472CF2AFFD02DDABFFF17782CDFCEA351C3847BDE52BD9CD4146D44CE623026950DB4E5B72F971DD8785D522290F938BAEEEFFC1CA6A6362A334EC95134AE0DDD7091271C8E0E00D6719484CBCF57536712D154DED7C6748C6217CA33CAC94D9C3BAD9FB13571DF8C3992A24E6063B9EDAEF439002414F710635B0BD261A7482ADD40CA74D3591DC12621B8BC706FF0492F80F60131A241739399D37D27CFCCBEE3ED13144EBFA5F832382669E81E3B68AB28C72279C859A1B8A1377828041DF4B8327C4DE1E0C9B3CFB648D2382712A8F011B564A806CDE1BA38F40A1CDE2D1C2E9BD5C409D76B25F77CC30A7D40AD645E8795984668E938EBA7E18934ECC20F4DAE563F33E76BFC1021A29A94371F57AD9336E967893DDCF293466255DAF00181BBAD785C6E081D8F3CD3CCF26E05EF7A9A9B367E48320B789F34334F5346ED6023F49D5CA008C2B8C866E09294F1880383CAE38EC563D690B34493544FBB80D5F7B361DEBF33D722D9D963015050F88F4554F7593A85F1E1AAC5C4FB4AEEE8DDDBC318F89DB31690434575ED8D6018BDCAC68BBB10610FA25B8E3CE7521911FC46D028323801F1A2ECB12BA7C3673F07769660CB4ED72A1B6801616A71C7321C06A0637F3D3A3DC3045A790446C53F4E1E85A3A93130D21C60BAE6B62F933784D10E0DB6D7772DBC0EB91CF0D7D90D0768F76709DEF4DC8577F9414A372EE8AE202BC886D8555486E8989B5C5F27B41F9E098CB829F73C97E33C22A431435595EC673EEA7EE6649828C48F2A78A063614227A4C4762AC1BA378235A785904319DF31FDC62C1A4D9CC60A14806F78ECA87442740EF365AECA36CB494541D4C39C5CEDE32690758E67561D8DD1B001BB1322CC0EFF5F45DBD62E8DAB75DA6EED8CB237F06F7FB3872DB6AD28EBD9245BA2E40C4328D88DE37910F4F8CF33CC176831D0972AC61726EC0766E3933A4171DAFEE475CF24FEEAF2C2F10874005428C03CEB1C8AD145133172DF53049A0BEF592AF8353814591BE9EA9CE693092F1CC6D99987EE4A9C688DA04E01B1BCA158341FACFD9EBF94AD5207A6EAB74B51500D8A2FF7DDC7B806994605F994FD1BCA410E4E67E8E3143A51D39A13C5F761587755A870DA14EFEC3C600747DAD49E7121BB7585EA9AE8E25A58150E8BB7288F349A4F637EE9DD6EDA296834192C8C4E5DA50756FB3C0F399B57F117171000831A7DD592883A31583760AFFAF907E25F51026E7EE89EA83C05A8C4DF9C1FBEA4C9FDE72E882E76C955B82E33CC78BFBDCDC3295F860D5BAA2BB454581B08447EE2AC774DFEC4042608C3100EE07BE69785931E4C6332918532421ED2B94D6410E9ACEA948F113FB221273E668E3163A1DD3DC1833F25088EEBAE3A280DB98AF0BD095557297897810B86B81297864385D4D0CD19765295B435018504BB387F58278A991C80DCB69F80CBD06D5D18CC440E569368A095359583A04A82ADA4665EC3EC7F5A8938F26D90BD8E6A29FAD8CABE532D011B9DA5ECEB4C9FEB6FF954893A00704CA8DD1B9B737B059685C31008C281EFC161DCD5279F90AA753F901970F41B5DCA7BD8CB90F1618BAD0B5813C76AB12ADFCCE91FFA59E5B6D37E2D39DBF4CE462DE4A4EB1A4CEBD239583F8BF2F6ADE1A37D47EEFA275837E9ADB7BC312D655DD628E857D6180A3E648661E479191CF6FCA305D643F3C1B62BEBDD8BB06271DB75D71B36D7EAE0DEA72549F1F26673FD566DE3CF80DAAFD90796D6C55E07DD22A08AC33F5B6C4222A2369B6D7A0D6F37F808DD5D4E2DE3CDD41E334F2D3F8C4D5853C19E4A2534C7EDD7F41ACC88DA0DC94513D6EE53209A2D53B10481563F49121F43758A470C44563A57B401830D2572EDA322655588713E92802DCF684A36EA7F4A0612A573618B3BBDDF23EDF345539761AD2FC779C2DC123F500D65E710F2331387D8F98118A5B67E92233CBBA0938572A01D17F8D524DDD99E62A92EABE67D1CE4B13BED634148A533C511302737E9D06E225B6468566A761D0952A2B22D1059C7D0A0F4C6113960D885290EC64C88F038A9445AE10ED0FAF804D69996690A70B1355361081C9C663F9315E7CF7127B8B0FDD013C9DA5DA61BBE565C870E6328B8025D8CF0C26693F5CE9105BA509934D3EA06F3C21738F68FA99E3282DED1B1CD9F5F24A98014A4DFEDD2B902AFA5003DCE3813C6640C6753E9F33B61297804403374AAEC9E0163A8DB2EC279DCB5C8A285A40B1FF66F2A62B4B8CD790F36CBD7B6854AC11D3C20E3CE2AAB8A36E04CD3DCED225B38F30486A8FDD79C40EF2583103AD20D3DCE0C4561D51A412AB5411C05F444E3A613F7CEB6806224987B5FCEAC4C0AB0043A22D5AB7C6F1020CE821FB302E0FF0F3F5F5DFDEE011822A313DDF94417E84030D74DB9696B7E192BC35E35E620D8A26359D1FDCEB91FD3096ED8D91B17C4854DD6459594B4161EFCC5804DA58B98E993828CE597BD6DCA010F70468054829923D15D0A1A2250BF58A3D062ED34768495E166B3FF18A59A01E25C623326C44963C17C79C425F9327C59F4249F44D3E2CFE084357883A0D7007DD188E4965E13C1CDA8C9EC77DC451B70DC91ADA52EA63DE58E7760524D149C643D9A828914EBF1B121302F243A9F3C5B2718A0986A4D2718B31E698FB329644A7C8D5FE1C009C678737650B2E314D4B64BBC4F90D4BDE0EF3E1799E554C908E074A6DE1CA5112091DBAA830420612CC518021A074DA4B78402CC052E07B6FDAD67289928F6718D31420AFD3D3FF83EE28539101990240C707277D82DD339CB00A4CD747C347F5FB71695AB6E79091C1C15A5D6FAF597C1EA09F3C4A55D23DE81FCC8ACDD4B2DF614722D18B9C5D89287E8E007301D3BB37ACC45F93D449124D2A0A75C920C58539852D5CAD778615FB6D106E159BC09E0769D8DF33DFF9CB85294C0CD847BBFB404AEF7F18159714F4AF9AE2D15DD30722EBC2D2B7494E9A022E2E15229DBFD06890F397ADEFAC18D5428EAAA31D0D1DF1A695BFF53D7BEF06EF8DE07F15ABDF4709A8096ACAB57663933134AF1E4ACACFF4CB98A3F61C8FEA26992C9950E6E10E03460351BAFCE660BB441E3419E32256B412E42831CCFE11F63A06AD39C66625C127AB08240D65EBE596ED20234B64463F6E0733BF945C9329C92E411D22F3BB07FE34CFD20023C74F21D9797DD9053064BE94206628130478385A7D4903A74CD1358FDE33A74807E76F27C3129691A6D9FD3CCBFBD5F1E3279964F6701D83E757F5865A14B020A62895F3FF8B2C57297333DDD5D74DCCE31960914828BE6B3ADD5D62430027932A2F35600801BE105F1984703E22BC961617B91AFAE08F815CC8B7F6AED9C55451DAB1D3BFCBBAD6D0A1C140F5348E971EE0EC8D27D09126662C3571D31D7612BBFBD8E33BD7467BB82969E6F79C9B23B3B827D94ED39CBD27600CB173A8C29A5B88AB661AC929F53060F2F5418B42DC50B9621F788497CE0C93E4856BEE0B9D152B55FCF9B434CD2E916D384835FCD3CFFCF08EFC4C54DA50B68089E5F23FDC00483A67C6D302F1AC45E162677F4EE2C233C49F08DC5B276E4F15ACAC032647FDAC14C1EEE18C4A95849F2F96038727D21E1258AF2D796022E10E8783533AB5D19C4BDE7200C3AF882BEE759B66E5F58A975EE63F62C5ECE3FF15BC8CEFC5D7E0B3DBF30939C0709AA7C48FBF2481597CB8BDFC0ED192E4471072A283E2D9397B6E44F23CB1BC9BA0F4FEB167D0F12A0EDC8B92E4D4069A448FD6E122FA7D6FDF2B1E139839EE31C788E80104C67DFD3CAB321EE561DFB5820DC41CC58502A400AB78E017D03CC129B97394D33B1D7FE2008D691F2ABD24D7CEE2EF9A244D3C8B6A9070BBB507545268C1B938AA48F8C0808ED520FCD761AE837A27262BD61DD5AF07D302FB6EDC5E8338589DB0E09C3B9ACF32DBE317B1007624C2C70505B0F42A8C780806BA276392D4B49ECE6DB836587FD208410F9B03525E6B431D8DB0C0D337E2EB8984AEE0A917AE35C690D6C24AA2465031BD1EF28963B2964A97B2E0813C880FF4A8E382DD4C0146609A195AA64DBBBAD81604D8B11FBC02468BD59A85EA91CAEAAAD4F6128F8CD0B458E11B0A2E2BAAE78A6B23E63C543EA1B0CB69CED38756EEC5BBE89392F4A9B26970C51EDDF23D9D32F434D876A0B2C7BA91456A21547CEBCFCBF056B90F48F01994311704664D197E60AA564DA81C5B8AD70EE289EBAACF37CD9AF9D23B872118E92ABF7D162ED1F5BB2348203DEA958D1180ABC6756B318844F0924B32203D0E0382AA1D81C749E4D6048CFCCF4EC259A9190D716AB29707A8B012C6C064B894D2FEFA5561C37BE19BF419BC88C82AFD53E649A6C6DE00B233CC9A31AE4A0F619F9E2C72B407781C75AD02BE182B0EAB2A7544245331368DB373DAEAAFC4F88FB3E2543AE681261F6E17E32F3DE7DB31543219F1D79E6EA49CBAFE608ABE0943C8114420781EC1F5F9E0B9C94FB08561B8376E7DE8846355DE74C1F3286FF7466B7F16463D10DE9654C424BBE8836732C150F810BA9A8BC110FDCFD959CCAFB23C6333A39CBCBCBA6FCAD5C9A67AA00F92E499F90279AA302F1A0D7E9643D3599CB4DF568CDBCB4FEFCD797984EFC9232D18F11F9A67D16B2F9E79E2B7F8A728F95593CB98A1AD73D62133FB028EC8C648F895EA9077385ACC647881D52EB00E14AC7D73D13AA4AA544C0AC9C901FD4B8C39A9E3B19BAF1F376E43ED5DDE8B681EDF7FA891A57BBA6B6E4610C48D3EFB549C801AD09F86E013B70EB7259CEEC573C219E828AEBA65661ACB5016B747F3865A6C51853C091B53D5485980EACC2920E6CAF918BA70168AC6C4FB0C6E1B84C79DED74B310CED201BBDE001DD23B581BD4EBCBD836D35F9CB43B97B56CC36211D9C11660B6BF35A76D35CCB2E3BAFB55DD56E608FACF26C4E79172B78BA9F41BDA3712929AB14D4546B258E1F2A83B7E7123D1BDFBF5305F7FA731ECA45D3542819B293EB9AA8509CFC0142E1E9A49A56DA58A155D8FF971160C8452B19CA1FBA59AE68754098B4D625535A61ADAE197C678E12F2A3955AAA6A28B06961AFA7F627F53E157C01265BEEDDAA1D0007E9898C0F1ED4EF7F87CBACCD4637D4C58B5A3367BB3E3F159F8B7BF7E6646DA93C5BB37986943C6E8900EE344DBF5F7066D7972BBCE7B80FD58425D0F05DA36AFBD3E551FA678686DF56FF9BA564A0FDBCFB72042B4A1C581946EB95BA020A8E6A55AB610838976BF3ED1BC477D20740D679E7EC62E390652900328F2DC75713ADBB01544B8AC68EF0E3F499E0820562FD67BDC9BDE1F8ABA63982BFC5712D71B0534BB525E4251E4FB907775688F360072352824491B9884BCA060651DC9C9BDC34BBA774815E4EB0117AD584E5DFBB74B837543199258DE5D3414724F99E7BE47C94B19E61E2578B01012C734F2BF2829A0ED375D0C1D74D74DE20147A0577F82E667DC42F7AA1AB794E94EBDFBCAF4D103C56774ACEFA383F75181BCD98DAF566C522814DAF6734125C8037E45F101847E8BA3C9668C45D8E82D4D2FF2140CCC0E1D26ABE7DD15C47CD98BF08FEB97D8AD3CEF63F0C4BF7493D16E3BF1485480B62B42BD8F7D51EC6A5B8C83036746D399F607CCAE7EDE14DC166CB22E53EEB3983B7154460722D4601C0E05C6D9264BF45A8390E37385B9CE1B2B565DD528EB693A932B24C9A0B464EAE56DA411E88E619236F7311AAB2D1B41C3D1CF8EA153FE134B6652A66A34DA0C456BABB313E8A287A2B4AFC4A8082F19CE4256ADD50DF4625969B5BFF89BDCB4334D577E03189A98EC8C87BFA1D53968AC9794E00A30CF25A7454F7DF3F99C683B910E28CDC0060CE7E12E429DBF70F8EA4DFF1152451068B37FBDEF14073DB7135A088949BA692139FF6A26FE0B5BA564422D47D869DCB18EE4353BDD719927D75880820A7FEF672532BFD69095340DAEE2E5FD8F899BCEC9EA320483361A0509BD1D4AC7F4C2DEE365CCF960EFD537FCDA4BC8D5B10EDFA72DDD56553249A89AFB590DC329D6A507BE8D863DB337702E66D214FCE4C965FE5E136B5BB375E37CE2787B5C71CE5EB65D539ADCCFB660A9D4232D690FDFE1C6D915B252DE10BE1D5121A10173F423F039E58E598B10F3FBC79300BCA7357E0741FBFEFEF149396B653D43DD12A8390608246C3C07EE45DF9207BDA8B1AFAC215BFE901324FD0FD942C3108B72084A93634315699B0DF845CF9311603CAB7D05F7CA3C68F576578E8A80505D93277B792F90D3EB5067764569520CFDDB6D2D3ACA895C922D9E329C40AF5EDBBEF7CF1C0AD0188F09E9B92BF081846B785738CEF4DF43363CAD744340E3959D1AA90467CC7A89FB8EC357C380201E00F41379BEF82B6CB27FAFA1197A8EFCEEA945BE41207305663C5E4454EF35EBD44259FB9C8367721FB78299CD418CBA9EC26D3CCB0879B376283A89C4170F03CE61690746FA292EA994C0E762B061425EACB8E990BB66D5EE004E5BE286562F121E4859AB3691145007200574EDC0D8571174A8D0DA378D386EA10C6297C6E0973B7250F4DA9F5316EA44C145DCC187630E8FD076BE140C88C05FBFC9F334959A64D47EA69A5E778A16EDB073CE540AAF7F389846AD0FDD96FF4146234D55C254FAADE2AA495B35CE5B2875086287F6E598D6015EDCCA90B923152BBFCF166AAE56FB69F3C0DC74C7128A971B63A8F0B2318649C601C4AFCCC44A7062962F656E836454E4030DCFC69EC81273102C59A3F1D222E99ED13D2BF61E577F29B73E8CA61A7C153E7E5A0F5E1E5C5A39A16268DE128277696D0011D9C9CB478973F88C282436E5B98F4B2D09BB08B070A51A9A645166F391B96E8FBE837B792BB8EF420A78601BDBEB048356D96789D9B18085279A05C93F35694DCEDD31438991ACB728116D86DB69A78DAADA2B6ADCE97D91A153528F563B9EB7901D94F10377B0BA6124E57180CDCA892BA7C2C0D09C0D7691E7DC4D17584A9C261BF1ABA05605A796CE038AAE23622D19678F523D79E17EC0113E39CF15BF27C0D94F6E5DD4F885D569943A39F50990825A793F6E0A57A9C50DF004DEB09758044EA51214E6383110BA62B6CC50C8C2AA024917B8C9F49F946F86016EC18AE171975477460531AC31735D7DF7614623E7DF77EE10EB34A14EDF2BB910A8B892C7C4FFF5DAD418A3294B305C9F7C6BC108479EE2828957D30E8AA2788998BF5350A89C23D97FAA62AF1A2B6A208E560965425C308ADFB1481897EB0C851D54E9D5E4245F6AB7FEDEC3ED08CE005AFA59FCBB47DABB4D8DFBFA8982CAE49147C2340F8405E4D521A3D6C55A6B2AAA22571E566DEF117432E650FDDC7C64830327BF1BB07E6BF64BE4BC5DB08547F2F5A55BF47B317EC09DD481F3580039E2830DB6AFC87EC7DF6F61277788AF1D11E08D4EDE85E2EB962F6721C73EC75F8FF1EE7C5A35831FC87627ED71B27FA98D07AC9A156E1CC3E188DC1CF943524AB466FC9345B65709D35F811C623D0CA469BD33E9F941279589E552AC3397933DD0D51D49EE115CDB472404D3D0D84FA1304B7048B02B61F664CE7524C81C16E89B624A25288A40508CDC9BB2B106E03346CD048F24417B8AC2153579F9FA1511B447B7BDDCC0E8A4AFD5CE21B08529BD7074649D6EA25C45D4833C2327083EC0D8D21A296F4622B5E16ED19D0E93131635D8E100DE05A213F309D4F67B68859ACB069BA507E438217C6E5A03D603DE8E9A737EA0CD985D014A8AB7CCA679935D708D5AFCEE19585C631D78514DD4F94374A56E6514D8720B08684E68154813425003F047CC97F419F680453F3DA090B21E8A0DB8B78343FD8375C1E44D27434232F0D38C1232DB10182D0FCAAFAC69D5C510599E3F7DDA99095B3BB3D71B96F274A88A889D2BE5671F377185C7B95B7E09955314BA9C52147595E289CC8D0D42D06D894E13A4077154A0DDA0EC4D5BB76C4AEF1676CD101B1873C36D9516E900273FA4768892A5E93E116D0A90251DED8805245EF3111D3C462E32C0FB9E329BED9D21CB8348962BCF8E72950DC84531056FA4D260328F4D7B1C11F5AAC696AD2D3D34135B3E3E2441791138A058AED7B094A981D020F4F246CB005F26F664896B4BE0C63C18FF1B9C53D102D45EB55A02F414C96DF7C6D5D866A19057C5A183F69987D26FD111DD0B6FFF3FC3CE46FC307FE40774CBA58982B2BB624FED8A64AC2693261537B9D379634317BE5ACF0A4A3977123DB9377A483C73C04E5654BEACD67E892808F51C30E75825B987B8E6852B741A9CBBED9642D208F7244D8214CB9E8F742FF4AE343885B3BFAB4D20B9C992FF0635F8B06498BD41A64326A4CE59493D5828F759E58E3A674C59F62E837F01F0FA6201355BA2A09B1851925A66D0264F251E01D1906ED6D146DB1C6516A88D941DC358031B0FAE9E7FB6D808032F67F4FD1390B2FAE2961EEC51932952A3C0FFEEB8ACD7E29950A76C2321175EF4AD8CAD7A3B69B6032AE21D94FA7552C635791D1D59AFE8DC4238061DB29453196EB8B7D794C80CDB7334D47FB8B66D2E21827FA4E04A24B7C81C42B62839594F4B5ED96D31ACB3FF16499E3A630B7446D461508A857E44FC0E90AA15FBF9BFF5743B88EF4E5174820C9CFD497B69375BF7F8BEEF4C089E3EBF0211B943FF6ED53D73022710320A5B06E6C264393F3917F70CBE848562501EDE7D8B3BCA14BB19E07A3480CD3264265C7001C3B1B7179180A377CB58730E79564F12F5D10182FC1EC632BDCED37C5EE67DE925D67430C28FA18ABFC2E7003215E4561A4FB3880D41BC5D7CA583D5C960402CE2F6B2518E2C103B53E2CFF94E804F6D47F72476256E2680CA685EF536BA7DBCD2013BA561EE261A8DA559765A7D57AABAC94E3D1FA1B1316A8F56EFDA81FD1657EA358762FE7F363D31BFD52BC74E730BD0A177115CF9625F2277E6242A38AD92554507CF402FECC017A7E9937407F25ED06C3A306D1D268825C169BE2ABD62291A260CE91125D42F443F96710A3F4CA55BECC0F74BEC44D80DD75B6E982B12660E6CC1C7FC3AE1156EF26D32079E68DE565141671571125FA6C00BD9B74B9B80309D2991463E794C8FCADA074DD0071E9BBD8A80DC953744012AAAB3E2D58EC0C3EB7FD46C5E052BF8A12E86E4F8347A7004C963F2DEE16FFBA71633F3554F1C2E3CBF71DD1F2584A38BD7E7D037FE73EDAF3DB5ABD292F93C0C1A816B99B133A2A7EE8E43409E917C8EA278DF7AFFB88840173E2A7DF81A06EAB17BC1853F42C96D0255B950A54CED71B3CD3153D159B0CDD1706DD4C4635C9F0C71ACA9C43BBA22BA977E4EE74B3630651E27EC8DE45B23A31BBEB23E6B762D9791EB185ABF2E4E908376EF38FF65E5EC811BA4AC45DDE55E9E39E79205C73332AE76161D0A0B785142D48FAA295E65E142A24760CDCBB4F5826948D32CC6C74AAE369B021289C5CCC2AE81933C8F22549620C7A513B07B0BC4CEDC52B502DACCC2C4280DBB04E37C13F4E005CF2659FB9957AE38BC2EB0A2A0E8FD25E1DC90BF582E1E08137FDC3A28AD8B3872FFBE55350C85549669AAE7F1A03A66FD2AB40C8F06911FC3B1F287BBE3E26A732F5B533F4F377EBAA2163ED895FBA49748A2AAFB3B1E5FA39B9E959E8F911A21E51FBBA87CFE01ADCF8440AB7BFF5AE73D625B8036DE0A159CA28BF4A0212016ED0629DE75C8F9568DE7B85CB5028EC0870E755F364C434EC34D165DA712AB6185B07DDBE1DAE99EA89C0589CB1673865906A4711584AD2BD9AF66B473AD6C41CECCE4FDDF222D8965C8996BEFAEA338D6E7CEC14617239060A6F9077BCA8C60726463F3BCB6DAB61FCC34B5A340E96F2256964B5EE5EF76E924B4615A4A370DBCBED2E016AB24D35582D7B4306DEF2718DF6C077C3AA45F53DD7A67FD8116207C63AB1D969F66C29CFE7C13F525F6B165954125985D0EE82A40BA8CE850E2111628D5744F4CB9362D98D94CFA942B32949EB0F55F7B3B27458F81C857DD7A66E933F409B575244185BAEDC29D3557F5E055D8F7E0F8D893480D276500A89FA20310032FF26CD6DD22DE2D87201CFE6E9D685A665654C4FD8B1ED49B2933F31404408264A2D3BA1DE73BB83853FCAD9D040ED18209F8DEC0E57842DAA3BD063D12DD1013044B8A4ECC0E6B0469820BF67986D461A7B3B905FEEBAE7EEE51AABEBEAFC4F51AD370FDE1D67F5130D46E25D9DEB2AD2A2CE2D51F73A4A7E50F051080C5AB319D741C7201C75AE181BBE457B49EBAB45D561A5C053EC9D21B5C8BADC424E15A116A8060042B32D1ECACA7EA477149BF4E2C7331BA90E80DD8CC2986FDDAA34DDCD8289D95912908151623E75709BBA7E7C8D69648D3A4B94081B243C06553B0C699882C85AB62B1D27170055FCE802FE9667D134FE262A72BC05B5FDCACC01C450D5B44CBED9BEFB7360FFD352D997B8AE146ACE36062A4DEF608A5BF735276A1C8B8F2252F533797C7E45ADC2653B8096C918C87EE8E0E3A1CDC9D9F3017EBA8CAB58B394A528F9F9B73F6158649A9A09E4BAF7EA2E289F50AFF86216EE954D672215A22D17F1F253EBBB00868AE0A3146E40A0E6FB8E59327B286DA5AE4F459CEE9C5B947A4176A8C5A3F64BCBADBD133F15A7BA3F62440DF8A67B785026199022D84CF01DA717E23C5418CDE5F7D4CEAAD03CE42A0B64803EB6900A10F4B3B107A28249E2413C24B0D494EB2EB043E0C827C025D27B022286ABFA9245D6895B6CC4095B7ECB4380ABC32EB71A649F14E047BCC6174FE7C323D1DF15B97B4DFA5A56265836EAE3AB06E2EC2591090E2AD3E577751B1500553FF6135EBAD6B986A09E61D5ABA190FB43AD5704755F1439FFB113FDAEEEC9128A4FFFFF22CCC650D52B174AC50BEE1AF046E534246E150AD71438072D8B456C12D6DC6DA13DEEECD94909675B7253A3199EA3AA453AFEE244DB1E98A922D126FCE6A86BE7314C08F4B3574D51EBC800257E7A0AA04EE5F99BD1E7977C3EC43FB2B4599A381851B76759592209940CD778CC5DD55E082F9EB8631DFD2FFC3DB3C2687A30BE6290978FB4EB94CCABBCF274E0BD28EF172334931D0CC9B815C2A6AE735900A3253BB70A148EC3188849159FAA084DB0089A1A40648AF318525EA46E3ED1BAD118B1D15B4F4F74EEF9058FF8C65C5FD3C55A9705A87A619160D4DAE9FED63DE72FB19B11B2E09FD431FBF47D53045BE16560532228EB14DEB065516B3518CE335647557F9D4A872FB2022BAEB5A0718E4FCA33D5DD7AD82049326FD0CD31A998F2A71A6460F646DF02E9C774FFC74EE12BFFF06D5A5DDF10A448749E20E4521D81FCB46CB7C93E54C350B8B74F58D640289DECA8C905048A6E5D71622018EB49A38F7BEB1735460BCCC3C0BF638DC91701A453625501889BBC13C897122AD03E3F2E2AD7814A8DC7ACFD8CC1B6C83D95CD626381DE3039A5A62DAD07E31F272D523CB9A6C6574FEDCE69E5164090FFF865AAB8BAAE934535B4B356D485B82031D00E75283CD09EB296BB4C4BD858B865DBC420800B960C1C64A3B8715AF030BD4423E6783F4B93B6E4E2D677DC809D146AF24BE579167B19D2A3C75855B36AD3B089E2B7182D328234321C5C12F56FEF2D7FED958E32D47C58969780AD887127FFEE9E42B82BF24A192F1B47E16CC82FA5E877BE8F75EA783DD871091C0045279E647C71956B63E1FB4CD13E9DAE0F5378A2304FCBCFD016A697004223CBA696F1C58B9BBDDEBAADC5D7C69790ADC9BA1F173C1BC8B2032266BCA019EB9F0B0884E68F3513410C53FFE1B790B4907AD1EA9AFD0E5DA923233170C96D01973C4D587644A30C60720CE7CC81A8DEF43702904C5907AECF788C4848CD6E52FAE9B1BE5966830F101AED158BE492F9CBAC6CD9F3BE400B7F4358CF9529B445FA2984A1580FA2EB8C22DE572B9D02F6B5584FDEC725A96B345DCE4693ADA9600B396CED6BC17ECB3C80DAA05AF669FE1FA5D8B9643E2210EFDD4C54EBF4A1AEF65D43EC2275F1752056A254FC28A3719F7A35EC77DEF17C687E8A0F684784CA44827B0397CF38CFBEA201CF0FC17D02193510D2F5DB3749F423EDB9CF2E7E15CF7F4C9602AF3F2B1E7D3A933E8AF1218B80510ABC4A21E348194C020149D59A0B90AB765BB4301C1B0600FA97A23A61C58F66F9A818477E9079056E7C72CE1921EBE807961FB5A11525CBB312DD701074493D10E40D5E7846555C377A21A2A92D6B94B7B6C7EF06CB7243BCDA35BD83921F8E8F54077DF68966C7DF0DC8DC510B910B1CE413E64EE5E8A7DCEAEF9D20B6F8D7E608D9FDFCF46F80AB3D96F3B901233B126E77C4F7D687029BBC7E1D9062AC6EE558173AF50F7B84D7D3D36CA808C8652C316DFDE021A51BE08A995445067EE51571D47B360622B5B5C3C7B7FE9E254B587D5375CEDA31EE8FD1A496F60002AE444C729D2E8BD286B62A7D0BC43E91BE5713B88C9512721953C61E1DA0B87D469DAAD2AF7E6AE21C2391E150D5DA364AD3EA46ABFD34CB24F2E2B91B8E94FAF99C0F20C1DF6FD81FF028B6D04FBE0EED84CD7F8CED0984112A884810495C11548AEB859608AE90553112CDFA0CFECEFC7B392272694E206D0BB078AA554A1B1C9327C30E6256EA377F2869E775BF131B2D8F50CE60522FB0942D532892AFB078BC1CCC3C6607DF37A1DBFCE78E92ADE275986630583870A9EEB86B658AC371FF39EA83C25F510E52DE5ED5D0C031481AF13DCD2F3BD15BD29D5084F65C175C050A7647560F6169A489469B047FD370ACBB6BFF34C896BBAF82B5F032EBF5EBEEB4E25F4EE704967081A43510B186E35693593D5B0904F51FF885FB3FC5940523A64CD0BDAAFE13C6DEB26F1C539BF15A672B56961E41195464FFBE7B898E4A0B0818D33319994BBE972A792F8C208742AB042E2452182862CDF7578EA78D52ABA0BAAD79774F51E6F7265CD5C38CA2926CAC62BDC6FF1741F2E36FE552645CB3683F9A7D2DC12BFD8A15F9346B3047B2E14B513A6D1934013338200425E947F8011323C559072FD9EB838E263BA075B1D207AECF29B53BB5A490F7A31C5992E21856771654EAE0705D9FCECD866C384001ADE166EFB028190F087D17C29AA87D1EC14A3ADEB40B1B076548502B9DD942405D93C01FDCE562AC6DE673EB6798F333CBB8B110A0579BFE0B93AB6B927813E054C785393FBF10E32D557C26697F50EEB850E0BC52FF977494B21554782BD96D341C469AA9ADF9258A74C6E0C0A0F9E71BC09532848426CCE1682342D7C8CB3F4D509ABC7B145E6CD51FEB0F06A0F2AFD53173CADB5D11EB44187A59ACBCBAC953766758D99977996FF685C0E5F69A4AA3333CF9AB7D97C62A6869B4E6BBE6C7D204B78392DC8BCE9ADD8ADB3AC6B0752E153043427B44D154E5E2C879A38F1ED0CC2A500203B976EF303D8A432235BEC8E117943FB882D90FC346B1658E954767772C68FA55B58A7B463BD6281543A7E7444F0FDD4140D5FD8C78A1EA9C99F27762D108ED4EFE91E4DD269D9AF01138BFF6EA6AECBB80FE23287E2AA3E6298867ED88283748E21DB6E3C123662649E124023CF6CF7902BDB03935FC496BCC5B4E5948BA167BD7C2589CEC444D37594EE9E05F032AFCF2205F2F1B6DC2126F2AE499292FB8F97E4C61ADAFF16904296BA78F584CE30210663C25C83475F399899F0DCEC73FE7CCD3F2D5656018ECC491CD5DFB0619029EC8CFF95A13C38AC7172135E0034DB24D59FB6EF57612ADAE2C66C0F634E500EE5C1938E987C57E8D124742A333F48EBED00596229805AEAE38480451F3827E3DE1FFA5E6B562FFCBCEAB6B6666502851C9D162787B235687433A567434D61DD1921A0C5FC6B46A9728FF850B74C856A3046BA5E4050ED893DD7B5E7C8EA9A5DC2344D2D3BFE93419C2A3F6D1E761C3F3E9E0EFE16838694D57EC3D5F9027542163C69A537C8A92D602D21CCA1246C0D03B1E549551C93D70DF28C4240A180023179CA7137F4F4403EF7F0692804D78F68BCF3C536E781F4281E3AC276A06747A0004E2F3CEA8F79D5DB17DEE0BC632C95F39B7374C988398EAC6D7F648F2CCCDDCFBF9C2D46A520645C6D60A775C3B423C8AA6CF367A4E0578A3D91D1AE8A13A9C69B960437DB8114E125478068F37BCEF4AC48FB5A06CB5715ADD19C6F3C4EB90998A77E492F1D56202CEAABA96A5D9CD6AC06A1A4535E294EF4BFC3C1116C3FA16496DF058F841C9D87A04F79EB6E25467584F5B1E002BF31BB2FE2F407701E2EC7483F0E23B788ECB6E48FAA1E6B49A729D56375D0DF8926334308C547386C6290C2768AF0A8AAA5D3689917A9A59BE4517F7B988E670ED5F85266F82FF76E3506814532D8F867008714A038CE776F7E2B8C9A4C148C7E8E7BC4CC45FDA27A0A5BC114FCF88832B28C044A41D70327532858976739D8283F2D7D7ADF706D7777B57AC5A12574F34380898B85F1112CD5530FF0DD3A6CFE130E0B184F91AD20F605AB41CEA344811E5606BBD787A2BD323CDB70AC408DC7A3D92A429A4CBE879065AC01D773F7B678193D21E5B4049977148594C8A909FC8E272F1281DD24386C518E694E9D1BA3297D7A2C07249275D743B46512DB3A12602BF5DB3CD7C8F113BF7590EC234801823FB62658E092D3050997370BBE057EA30FA50C075F6A5D8A6337D5E4D3B7DAA516C37CC166A150F98C089BB7D54527CD19C9D18459895EDE82725B1D65862B1E3363A0D9A3DA7DE740EF0E699EEE6180A709286C268E8EC6D80412F7EBD53A50B92959D43571AE562069C908DCCFAA491CB5162E553CC2E9EBF46C6124E9EA254A71F1A5E168712906D7AB550BF2B6CB6D60E04C8F2392A0CC9BB980212DB515CDF7100E457C0E4DD3AC8FC939E5E3A426FB88AFE7334007A401C835BC96E838264D0BA8AACA783CDF8767B74C99EE590C3CBD0AA605FBCE8EB93E9F5BB9B184D9EE8C6E5E0BF8C00D39EA6CB9D8984D6B01669218BC62347FB9B15C9970B847C9A08008EC3FC329C7282E67C44ED844856AA8A8A80B2E7D81C9AE6607C3F61EBCE95A5438470AFE70D609053C5BB0D4D65934A73600F248D4C2BD56D4F5DC6AAF00580F9DBCEFB2BCDD7C11098148FC5EA829AF38F480424E57542C376DD49D6813E1F0740BA90AEFAEF590C855EB878B505B70025089896C4D251DCF7464F187CF8C0A3D6EF605D8888E7947C4038856C576322B2BA1CF3E90035B88EAE2469FEA2D36456FD1FAE1ECD89932080EC50CCC6062EBC9328041FD8C08F235CC5DD24EBF237947D46E0C6E34BBAD76F71C748053600D08871AC266667A46DC4AB10741A9CB92846584200E497A51A59E03E06CFF5BA68DEF19A05C954AA807DB4C82E4F6BA8FCFE59F1252740828E030DA9E441511F2A78B13D3619AC9AEEFEFA20257F59FF0DFA06005645F0B7FF1C9FBBC99F39A13A3755841A7CF70F39CFC0087954C1A7ED0E36388628038DAE4C2D256EC7E84FA4A32061AA1CD04AF0DD003E99A0FDA1DDE3055C2192CB052E92CB9BBB13808A405CB50D1BFEBE3EE1FA38F9E91889FF2B82DD3CD2D2CF2F374A414C26A20F72A4805A9590977043F854A876518168AF69F43B2A01BF870739D23B9EEF5720F551C0AF918BE9B22A400E7E720660BE200B50ABF2FDC4EB57BD7C3A3067C0B744389469C571DF9D330B512263FD589B55BFFD44D1C407EAB6301CBB59986B0EA80FB146CB9FC7979E1CE8C86826DF3FBE314EA1250C6469AE84C55E1A9EC15AADCBEA4CE0AEB40CE6D2010D720B2F74B34C7DDF1115386635871DE19E60E1DE3B8FC43DC709970407454606066FF7064C07334C74A479484AD30476C64E6BBA91F8D9291FD198E9B2FB0C6A05C86F958F534CCFCE48EFEFEB56D0608D82462030A024B9D43A5919FE068B054E4FBC7A90DE9136A1F498C2F572ABB4A91665A971D527F19F11E4ACA0EBC72E03735DFA728C08D5D1BBDD53A0FAEC3A947F39FCBC4CE0BCED31CFD6E5DE960F10EC621B1CAD93F78B9A305A82F678EF4C2D5A6BC4D2D62C58066BCD3811235F1521397E9DD835E0C7D878E1FF96935B3FBB48ACD0283D47BDBB6CAB266EE23FFB1A81E7112C3F5E4E692F133FAF1531CE03E3C9AFB6BFE89B2824E7B3CA515D0FA9D4A74B354CFBD0AAE9BF3635D0A23441DB1F32A77DB4630134B7A81A6E33568DAE70F85701E5A920FFEF927463E16B60C58A211C82D1DDD448B0CF0F86553A37BB4A3F059A9F81492712260E37DE4D3678B58416B3EC07C364B1CF8BC3A033CB23235CAEBBA135278DF1FC368ED1E80EA6F017BE64FFD64CB265B70033A08F94DBDAAA700FDEB669E1FC1C6ACF93F7DEE2B0B31A43AD6DE01753A631593DBB2BAFEE41B9D5D318CC250DC5DEEB48EE4998C2C2320C2D3D8CA6E32F0F68112F42CFE1EC467DD7D90A0FF6E03008C628FFBA75B172454F35E63EC3ED5BE230A40E51740A85C91CDD0ABD44EEB057EBF08875B9590DA6081A70F1CEA241CFD24EE5B388F09FED5549B2FFE73D2E02C2E9DF0B1AB07A39424731F06539F7B210CB0889306A03B34ADAF4E84CBF22A0387802049EC2BCFC95514A560AF53781DB9061282BA662DA73895CE766AA190B6520D06720D8FC0FA8BF5A741194ADD6DF957C8C30D29E575B9FE5EE6EB024704F06CC4F1B2FDDD053B4F4464ACF6356E2C6E4EA41ABC4A12F7BC71AD362AF657D22EBCDB363C31B1773E5B8562BAF7CA187830F1B1AA20597FB8D8A0DC0CC6428CB577AAE8E9C17170283EA2689607B6AC6AC2661AF2580B21574C89B06947EFCCF4DB8870E5C3EB7ECC5FFD86B0B51E72F18610D32CB14831E9D787F7491B7AE593F4AD6F9B4181B2D2CD3CDA5C82B1FDD5594568D3197275975139902F5A5720643BCA23F542043735CC840BF5EACEC5C1189514DE081ECE6F06DE4D20042933395B3B45707514FA39C5009C78E28143C9F997E013BFC1DCF8E55F0B399EA4A62288852F33FC8C317DD864811E2B3D237719A5B8C33F6FDF00B06905F23D2F4E8836825F5ED81B0F69A366CDC5463889B391BDF67176E63870DF39C3C9DC2B0343BF69A2ECA2893A19F569FED8DD8FF264A10BB0426A6851B42D4668DFACCF60D2A7758A759D2E6813AE47CD91B2DE4053B2EA372C2E94303CD753563373FBAF747AC3E8A5068231C8CD227B811C3AA3A63D26FDE2A85D9A27908E18E9BC5AD961018F6363264C4B5AE4B846BB14629984CD78CB0C298072887271E5A81244C779D8725824BB8D3AC99B4586BC17BBE82F1E16689A860352E545A3816D1B2CDF22300D2C428ED618F6107E8395A2BFB44C8BA75ACEBF7F2718B84020EBB86945D465E7EDC610598693E44E00C0F11655675052FA1596C912E84A0D15018CA5E561EF58E2B6C48D7BADFD9D36A85A74E27E30E4DC7FA61DD5269E64C9215584915A0C599A7F211D7088BB7A00AD147C4E1AC9B0FDF4762E4623AFDF9037EADC3CA2405D82668F2E03C56DAE28447A66F94F7AD44333652673A8E55F2C167D998C1B921C6257ECD99D606622D1A6B7B06F1F2E7066FD2772D4C33DDC5C1A5FD9C1B960B58AC4A17E4BA79AAC58B8CA6966DAAF14D61B9B2E77E6610A0E4230E158483A04A851E8F1F63EAD0B8C26E3982F0598614BF1F202DD41B0DE21E44BC562E203031D71CBB7FC00A799F1B1C0AABEECFABA878F010EF5F34B964957BA18B52B0A5DE99804B52CED098603F655F3F4E383A631605F5D8987FCCD2D601D5879619B0CA49B55B4AFDF195574068C40A71D5B0215AF8ADBFEA03FA7976AF81BD7D5487E84789EA0A1B41A55C2E26611875D260BE02F4AF2E7A66D5312C9E561B6CB213BDCEED28AD7EA890C213DD92758CCA36836A77D5F1017C1AEFE1BC8DADC12D5ED64A7815A56F6A355CF9DD25B6DE370D4C9EA86F97913319B0FDF729729EF7C8693A69C6AC17C3EC8ADE0E530AC9F9733AC4CB6171239E113C8D7C7FADA46EBF87B203EF412919ECD5C03439A16255613AC3CC1A829990FCDC1369CEFE6A5C9BCD25F7B476364B9A969813B57E1CD1069F3CA4E959A7BF1718DCE971084ECC6B7A5C2889053F7EEBD990889BA1E15E6DE7A021140FFB264C4D32AB34F6CCA93C0103487438FE26313E5FC3A333D754F33F33BA588320AC7A4F3181CA2CF234E1B8A5B831E9AB5DAB35BC7B826E152F300481DB7FA74BB795188517B9B5EA86A91E5E9AAEE6C0B8E1A77A01506616B5A40CE7C67F88B5542F0EBA5E9D9E4365AAACB1CBEAD207A93A9CD339924FAD5E464969C0CB4C06D9B8DD9508CE44BDC8A4DDB2A7F9B30F5F6122D7B106DE342C3388154CA41CA612E77B59531C1112FD0999F641D6E165490B692F"
	// },
	skb := hex.decode('198276F1CAF3AE81992E53BF1EC51AB370E74A22E27CAAE9B0C953B2CDF36B04EE9E93E95DC14F02AF76FBBF312BCC5AD207561EA17CB649E4CB3FA0AF5F5C10')!
	pkb := hex.decode('EE9E93E95DC14F02AF76FBBF312BCC5AD207561EA17CB649E4CB3FA0AF5F5C10')!
	addrnd := hex.decode('201FFEE926EBA71B8222D98CB8CC6BCB')!
	msg := hex.decode('C09D602B21F3A0B10E4BAB37376E819F1E04783B8BDD4481FA9BE228B2B33F3686097B0B414C51CB51ACC480526CD8A23A91964B84567B3CA8A27873BEF15DD2CCFDA40F10BC31B54FFC920719ED23720FA11A10860B342B188BC77202A1C7E3B3DE6D75DFE74355A21C57B88194C870147A1586D511B0397283F65411D3D1A7B5149CE15D38EC2527EF223745A6AE0FE0D946D3497DF750BFCBADCC0C6B44C4539D5F30A4A8495B4E5E03CC617005204F03BF569825441545408AA6933B842ABC83A74AC7FE13A02FDEF98E923C904971410790960048FBE8272FB748783A47ED9509F2BA776157945556E0202D3C74F7D21FCD8271C0C57662C22955A8F685BF19BBCEB1881C900E8A0257C6BE5DAA50855F3FFEF961A964BA7AD70870E197AD1C9F7DD78DFA57121DC7E41A2580F039CA9A373FA3A25E97935CACDF2EAED66E1D7C46AE9674EBBC9FE2A158F93CC0665905B6474FB429634E144C78B7F6F4BE20DD57E6E74A3E80E187F4CD05ADACDFD463D5236CF64C74632DF9D5F5CD4493AFA705A51B95CA2F28233D9C288C9047E94145FB89A3652683737CB17A67A31F231C5A96F496201A5E5FC7D21CD0E7DFDE733D99EC67B0093DFA3C3CB0298FEFF55A6C106C6FBA26DA316239ADA220BFAF2CDA09579979902CC605AFBDFB4CC19974753D90970BB97C943265F7DDD042A9F938FCEB29646B97FCA7772837BB0D975A167DE5CAB9E728C632BC04118CD43D2EE67908E31CB0F25A08497E337FAF51377684B10D70907240E007D957C69F4625ABA8E60D450EDEC88B565A2B2808CD0C13CAB0D2FAE9D6CC864DF2FA787DB16274A73C4DBB64022757ABF6465DF88ED20252D47702BACDE7F5A27147353573829DB823B7DBD05EE842B38DC7D0CB6FF8952830EC004E1A985E171D1A4D45DAE572C712CCF024FA333ED5C61D532BFF12BCBE8D101BE64AAF8414DBD6039DBD08D0E1F3CFDD2BB723384BD24AFE9FAD3AED20B70A4DAAC66597F0F8A747337F101FC4BC0066ED3374C9DBBBE14CE19F7CBC230982ADDDCD8CE259BD11A080FEF32D1E2C9E1C695DF7A365E81B37A8BF540198284526AD2F4B62D86AC3E4D7D9B2F6F28A0B36A115E469302FDC2930654C1DA2E87932F4E6B829623F314EC627D342114B9DF5DCF6E9125B3A0D6558AEA20AB88A0CAB1CC342907FE82C8B273FA33D9535D7D26F04A7AE9396F6367737118FCA598D6A656878E91E0DF984A57DA85171849C6A3D6D6346F5721494AD609D796CD208D09115C231A0143FD34A9D21A72AA39715B07E61D3291F7F289A18FE5EE04421C725D2F508994DE99E408D65759BAEADABBE7EBD8E992EA3871D5C7E89B38061B012BC56D74F55936D0CFB01CDA79D8419A2B1DE41F434837BAA445E2DBAF599425A0D121FC74F5C9CC0B1C31DA94DCC7B89397F4DC2BCBD25DC1D27ABF2541FCF18AB1B73180E5222FEA1FDB25A6099D1F05081DAC5B2ED76802B2D1A725B3EBE641D7D431FBCCC0B1345FFB0323E510A389907301384ED95EE3A30E5196668FE5130F1AC6AD16BF881955EB348DBB0B0114780DA598FEE56C9E7148AB54DA072F8478BE2EF6251B87461C001DAB77D02C4E533B9D96045DD12E10EBB8ADF594196396AC5DE75964400593B9F6C0137D8A39E690E8F37AC630D6A5885A65212AF002C03118F21A12EF4C2F185C452476A66B50D9C8E5A6E994AFAE77FA48A07F2DEFFF2B46C9E8DB13BF869FDD1F65DF4EAFC10AE44F1AFF2E06FAF1DD2DC275DC0C27C224731677763518D3E4C4F09FA17B95CCCE7C7B45A2239E5D315F102C937B54DDAF175AE47C8F776F84CD12CC642C50FD5A65F130D9C6D97F578306FD94ADA0F79154BBF278E022BFAD551C8BA2F5E0384CB4DA3472F6226B19C3D49F4F24B4A148B5B254649DA2349A64270C31E3432C224612594EE9BD43B920901B14CD13C4614E6EE612127E6F1E292E2039DB8BA9EEF96C52F915EFB7ABC466E30CB05DB89450E7BD8D32158EA91B7F3EA1591810039CDB7285A82548FBFC1837A1177A8D67CF8941FB8F36CA6BE20B1E5EEBB3C40C17FA874DC5881D92D34CC3FC8170A429DE1A552D14380E1419380DC5B82C38C014B911CBA45B7224B656238D5AE3A3EFC0D68B2483D8C529C62B9937ACC3F906CA2EE035607500594EE905D961C44FB27FBA99B12302FEF4FE7230B4A4C10DBC2F8551AA96239A5A87AE3772DDB3ABF6D04E08BA80289C1BC976590ACF87F7765BD38D0DBB2FF0786519D9BF2EC87B477D004CAC37699FBC930CCA86AC0F74516D563B490B28F71CEA30141FD52F28940D050A43E954CC972C8836B24CDAB87929BEEE575C885C87442600F400BC44D9CF176154889E104BAD97D157B04B42EB3414CC2A08F7AB7E5982D1F9A07A3EFDEFF70D9FC5EC9DF5D8E74F07F6A60A162FB17E3FBA34C0CCA737311683F932FCAFC80DCA61729CA244865EC9C452A59A9955F2E366DEC5EDB16F02628EE27C37B1035A9C40A37C1294E51E7012723BB999CFF8F020E40FFA644E7DDD9521976306714BF00C3F6A925623C776D92A3C2F4CA794264572B8FD0366DBAB45D2466C5BE7AA5EA178612DE63E72E9E103613FF9B3BFDB9DE34AA0DFED786D5D50C0D90DB88A4A6A35D2FC832209802388EA8BD4390C06AB4414D62204847474E44FFFCEA672DB9F3568F5BA5B2FA2C97CB55461FD51AD408F7F7084197FD33B9D57A2C4C30CE8ED4C7925D64C961AC4A8EFA1D7B011DC9714C2CB8F5018086B4F425075E45BB92E9D1473C9E8B2035AFED0AC21DB128DEDDD97108C2B7601C0330E885FF119A545018CFA4DFFAA2E354EF70551E84B69C7A2419F9990CAAB8762736416E75251F432846D44EA303F6D20B146D70D6433A7157FB2431DD7D97ED1D47E3F075EE685CE02C61BE28F476494AD617A398D6BD0A26B65DDD82006F8A05FD42194D40A922B70546934E6028B4D8A6324D079CEA5F6030301F11206227C0B01E51A84EF07C241F4082361D3B57D66FFDE4282F3A234EEB673DBDCE41F8887CB189B7FE23D68B5A7D42C0394AC86EEEED5318EAA47139D64FCC257BD7A26100BC81E6A945C3C216CFCDA173FA9EB78DB99470A3F844FD9832FDC2E6EC5A271FB6BBD7025527835DF6102FA2096CD411B212D6FEC117BB93833CD0C821B927FE6FABE0CEB06A9F8F9331BAB4D881D403C6E39F145997CA9689886DF5B7168FB1C50824DE6F9AF5522630968CAD451CF13287DFB06AEC0693895069A5BDC6C029BE68F9F473068BA5930900602B54E6F22D2ABC77404D19BEFC97E5FB40885C2791C1E19438491CEEFF20FD83AB032B6E4BA92E19ED51EB9FFD313E8FF58AC6918DAB6456C3329C5B44AAC82BEC16F03A26DA85061AE9D2F517A5C7D4A56098C74CEA9A9B3E5149D0AF4803C0460344C405E3EF8E52127B2746A2A80D034BA4486A0F2E31DAF51E1669D71896111997C0B2CA1F4AA803D77B1B75915D67B2A8C8DF15D9DEC3F68F252E9891298D979CD8FF10BFAB14845D44EDF227691B4DAEFB00A62DAEF197D0717634CE0647C46D43DFACAA16ADA96E0DC4CB7693680559FD9ED9EDFADA7C84AA266D548291210F6485906F744A4CD4EEA0082A7641F6DFCBB760275728F3D34E21F46382970F16EE41B88A47D0105DC63116EDAECAA69E89EFEC92A710511C10D83F85A71306058EB7F51CE080CEB7490838A94503AC8EA79B76889D9ECDE45E980A16885A65FFDA5CF15B584D3A0078893075F4AFB51AEFC8DF0D12E16280124E691A804641797D2D59FA1E9B5686A98969FF1EE032C7B38B5DC9D3E32C335610F6AFD3E389E1894E55277768A64C91B3F03E14B99009FD3DFE0928CAC8D354D063C4E7E83A99C77EB8AFE93004B19585949CB68003BAD4DE970E7C516041FD3F577B193BD2264FA7BF187365E7954B7B5B880CC613AC4B7DFFB90E8A4087972B14D1C54F2CF00EA063C92D4F37D498A698BDD8F76C12101DCB462BE0C6B271EC68AA3A7F3CE338348079D923C917C32B9AD53DB17400D54E50013365248F193CEDF667FA00327CD56F4DF84261611FFEAB4F6FE0EF5EE3D0A43AB1B8B8A88179BB3A85E8166F7B0AB62C1057D07A8902BAEC0DA508D57673DF7D697B3C320180A5C8BDEA64D9EBB9F578B665D2C24E0EB5EEEBBA2826427824EAC2012870826C91E31A1E893EF1A5A636CC4A4E9A5EA27F92EBBF9F9363BFE74629567F91EFC2C304003064CDA1A1AD8A4D8CE629BF4D4041931832457191147FEC2BE09F30F3C3B3740EE89EE313AB1E051124783FD47109F5B085B3753713E8CF48E04CBFB39C720426FE315635F219CBA87D847AE3C8CD779F52CC66C8D9733F3FD4D62C77C682969F5B08A2E9A9477CEB7B4EAA5228A31E0CC486353211602EA01AFF7D6E0447F728D7A286E7DA3C2688FF772807135A3F514430BEBDAB6D41E1EF7C25CFD07B63A456BEAC67F5633D8243E19F53421D1D40CF4DEA68EB4DE6840A7B4B18BE6A699ECB6A25309A0E9F2F99AA0B91F14B5D3A95E439391A2E0F7CEE47769493D72D4F72919FA058B22508860597FACAD5CC8010DEEFECB9DC2F6A0A7DE2BF17263530A5D567BDCC6E1985D0F2154A991AF9D1078DBAC808D224D94E6B0E7137F5FB9C4F3014C4A6D30DCBA7F8BEDEB57ED519EF19B512C28561BA990D91D939C07D8FD1CBC86E33E9EBBDA07D4D698CBEE7E0454832B485CC67189F48AD9291AE49F5624B9C9D5E1A6121CE3BDF2A9D000246A0238882B6DFDB6D682789940AB9F880A8EB6A8F058703CDCAE894603AD04028DDB84C8A2EF1E1CCDAA12562E72C0A629B1AFADE29DFFEECADB67497ACB50F8E8A71C1151C949AA2CA936E0374B0833F804016495ECA9A9ECD681EC994AB6049A599136B6B8AA3B26459A9C37ECB55CC7F08420CFFB4279DDD2D9FC046FFFC7356EDCFC97D0347C24D15FE866877CB6C2965C8901FB7367563906FB34DF1C763DF123A4A387E32489961C4352A8B2E4CE0ECB10E62DB8591370847AF4BE024124B291196C4AC59DA742A6BA4486D7DAB3FBB947103128CF0A8FEF69158A67204060CA3A8366E08755EB421EFCB2E902D99A055BEE52B1FEED14704CC21B78F951937D3D89B174C957A7A9D22005E37ADCB1849E83B8C3CD9E53EBF820382EFFBD7214D03DC5B46E389914B2104042C90C9084F11B366B7663AAF34E1FBD526C59CA1272DEF01B61A29FD4FF3F37688191FBA572A488B9DFE4F3C0492756FE1D8843F988D1E4C4B2133979D516506A33F41A951DCADAB05352F45793A23E9B1C74FB4F996B6C9C3709705D64DC1CD44C877287B2737308C7ED64F57E1BCE32709E45E1EA9CF1A67BDD0880C3A29DB848627361E4AF296256D5DC8B01D8793F9A340FF2845536BFE95726EBD5C9EEA46876CDE75B68768080DA37215CDAFDA2B8DE4AA257062F1659DECA5B2FBA3C9E0739660F7B221DE4E656F8A36B808EB3A256A60267E5DDDE764919794D6CE7897DA2B1EB9E9FF96EE0B29834D4956F634807B80743BA30B914F4AF74910E978E9BDD48CAF3D6CB5A6DF9CC98AEE2D315CDAA77D4EB7356C67DA5B259FA6758AD4B3727A7AB2D1DBFEC938AAA70AE6EC75E99EBE9BBE2C5B374F3F80196B7FDE8943D471DBA21AFB99423B7A126DBBA65B74901E85FECEA9254E1C95AD6A1E3A444A1762B14261050823BD696751A954E5EDEB37A5C329A1A685B33DA7231E57ACA3CBBBC2A09347AC36E2AEA0742FD88BC4B8CCC2CADE0F06D90245890E3BEAD25DDE972A35199DBAAD0283D3307BA9CB3D4CE30DF1B58A3AF6F0DB3E4EF5AFB9B5DF1B1DFA15D8A8C6BE77551806F7B541937EBEF59FB178FB91400DC1647825579CD92730EA5EBB0AD9ACA32E86CC36FD9CA2C71A07568E074B0759D1E2817262A5DBE43CF551E35A99C54C2EB8C403EA11EF42D7DBCA3381151D82CDB955D025DB5CF289B648EDDE79A2E53AD7A424CDD51226B3A64EBE98659B84E3305CFD7E0024D3DD92D8FC38A3E9259A63981C9A00B329B6D3D149AE3A8462B38090C89E3C48D3F43F2580FFC8FA84F0FDF91CC84F0574F8FA39C7D318120213D8C53327D922937F606B9F75AB24EF9BA562C03D973A78B4B8A1C0CFC83360DE9A2C23B8952952BD36B403C7B92C9ABB098F0779F09D3FFB7DC9512BE0C934633358A145E0F92AACDBB1DAD736F67D0ACCA198FD9794373C7204B1C0D62E6F108C3ABE3637675DA28C9E0D28D9B2002E8A285950D9C19DF28FD9AC3D9BB74BE9DAB48A3725073226F172BE3486C6151F424C7821174AC41671E33D6A8D4E144BD394EEEFD2437B0249719A9ED80FD6CC433A8CB0031E7DC9A45C7AA10A7C978C1196435C93595ACFFC7C4094136873EC8447E625DB25E216F082482C12787E8A06AD074BFB5B142A6068D5E5356E4BEC888D1988069D3A18E23EB7A783BA37D26175035E55FC799ED0EDC3153EC455A829CCE74A4AE0FF090C5D4774F9E417237D14A98B1675B970D7646906A7467629B3B18C9BDEB4E70B001AD30F6C500239F46A5BB4ED0859B667C5FE32EB0023E06CB4C4FC1E0C8ED9C99793702B2136D6965407CA27E2DD77ADABA76D8DB1A2948AFF30A226998EFB348397CB8007620F328CE38D94AEE09C56EB95AD07C35C616314788D3069627AE29C78077F34624359AF30EA1205A8038D600B89137197AD8A1700E24ABBBE6376F5933DB16EFD6274A91F9F70E77863F7C248EECCD96F76D929757C96D6EC784EA0D18A699FC6D64ED76283E871D6009497B937330D044880FDDD77444C3AD72C071147E70CFBB0F97CFBD022F074B6A0BAC8D1AE187F60E8B9976550C0524AA885735C2877BB5D68674FB26DEC0118632D379796E25CA06339BEA3696418492E69BD2309D7E4D8525FB40AB9E39AA65C01C9690A81B365A87C340C4F0DBC1C72099507935E1A2C9641184A48051D98460EB026818A53C471508223047B196BA9FC0FD67BE1B50D284AF45D4524B52BA038886978661981DF11E9486B42778B9E5E6EFE30BDD0CF78298C9A0C33D55A98ED657C06B8CA18FB3F944CB02D37B4E500901B7F4E1805B48E22427E15C1735D9976A3F75D8B2F7AEE4D49C3855D9B6C0BB0CDA633F30E915CD991E74406488857D10EC8A4C095CE374E725DAA628E200A87855D4ACB2FA73F47B7F35A66C961AAF325147EA5F4900D1872629B4DD814CCEC4E0D67F27C7DE58C6E9850A3E6A9B10EAA83765B0C5895ED50C6481434ADE00796400F7A6F54769C6F8AFE897D5EDEBA77D0FBB91C632C5D87D747F21954176C21CE01C46328DFA53C92BE39B61DC498B962694C1A02D6980573A24EFAB22F2DC4B4A642F6971CE11C15BBF2FC32D12A2642A54882DB21C810F85C8009FBBBF784BA6B8747EBDA5EABEC273BCAE69161F4AC4AB6AAB4E8303CEE2DD1F5C7CD445086D98D94C5D670F84FFD6B0B5DB63DC95248D73F0B7D5E47004D1E5BD3ADA857339981245AB33C8389C2271230308A0C88A4A36F2578E907FEE748025AFABA770F9B3CE8C2C66DF5B8FDB7F5845C2F485078558E24B7F3708143EBC8A9F48040B7AC6E5F78DA84DE32C72719E86A4AE9AFF1F7DA3A72237EFBB4C247A5A0BDDF169F60CF45DE39475390004835EE24448B906866D497E0177CB43EB221D86E32105D070CAED67A1758CB721B8A9F323967E41F13D2CD3C1EAC0FA5C0F69112C5AB8AE768288B28AAA43A3311B58C2721743544349D1ABCF8C53098D7801F528CDC27A8B1C1A76FAB19BC2E8FC5024E45E726DF491DEFEC543BA90F97374267D3CAF91303D20E48537F62248A6EF8A1D5C7D019E7F21D85F02B7ABF09FBEE0D3D469D8867D81615010ED167A3E018CEFBB30B86457FAE705260EC1AE70F5625E60504A23DF354E04E1599966370E6DC4562CE5F21D41342E9DA7CBBB8642B9AA435D789BC5D30CA132C5B59C2974BCE1CA47F13AAFA5ABD8FC1006EBE670CA96E5C2DAF3E0281C475795A7B92A303E9483A23C50E9AF7D1E4168C3E22A5436DA7EDFCC581940940698DADA1CC3FD31CFF221301D5B4976B21AE434842EB52221A26BB66BF020C5C3BF879A5051880285ECF2974C85D946354BCC88DF14538E333B2B94C6732EB2897DB5F6917EB27E93C358D7BCE85D4D4732398AB2BA4389B6291912D02BD5DEB4BF8FA9C310786EC68F3312AE09B75C4DFBB0AC51D3720927891719ED88FDC6E5F6D17434AB48F7DE8B6E34B36B12CD32F69BCDE2BBD59623C4451C1856FA24B3F68DB0D6EA52E9C9A3583779A5CD7CA53F60D7ADB1CD63B7A85E878502AB36C2D7DA80D7C7FC93DE497FB02F9D4E825BDA2EC38DBD0C8E775588C38E2123495377C4C8281946C3F2FE84BA3044C9307BECB8B85C0EBE879FF2AA2E9BFF9252F3BFF4E8DDCA6F04827AC24C44AC81217414C3108426F94860A282972DD94EC53AC956C1663D554EFD3CDF55471F3A2299C7F7DAB4CD2C5A715B2623096C3161C0195B7ECF1AE97BFF87DDA0717AA386C59BF35F3B1EDE864825DC5FB944C6DAED40CFFA960FBE8D1732F9934374805DAADF77D0471EA29003F17E8DA800AEE92B2114F1D85E564D7C4A7DEDBEE277B6B38460583DF20BF242A848FC4D3AD79510A885CB2B33E21B37A5D24310F5385CEDBBB87F95CF91A0FC4035BA699DE34E9D8ED2F73F65727C040627CFA308427852A29A30796513F39FC530ADAFE6115F75755B536D9B0F87EC31D4B9B331762CEDD5908AFD58B3E8E240823EED6EADD8BFDAF11925205DE32D87892D4DF63412042E0C5DBED13A668E7083CB7E3D0F756F22AFE7537A4AEA335F5C27CF4259660BF07BFCD40D0B6FC24493701A813279AF587FA76C4012701AD05ABA30FCBB21F0AE4CB0B6BEDDDECA1C3765FA65CA8E198D148A645A1458B122ABB1EBC57BF9BA8DD5E51F5C06C3E2E3F17098D392B692368FACF675AFD6936C0CBD72B0B2CB8CC0498D1C6CC4993A0AF01420A7B4CDD02E629E80F8CA041AF241E3E530DED2F822184DA172D504D500A5B079BAC8D54FF1FE5193BAEDA51DEB0FF161A9A9DFCB69DEF97D04CFCE7006596EADD7EF1AE3A39D9F109A4CC71B95426141450B3E7F438858D5BC88DD810EEBD081F93A604C41466CD8292343C2A4A605D250DD5BD6DB67D8383B5C3A0065B833EE1F7BB19B24B21EA0D209E72BC09431E699434942D9EFFDBAD5950E5FF74EE2005F1466D68C9F259A1035C6D922BDCD49BC215F57C892F276524E2A5A4C2EE6A8D319D99DDDEE07E8AB01D5CC5650090FEF5A8EDDE7C51A28A234C49477C09BE6022D292BBDBC943AFF371CE2BB94AB16D2A22AE814E8D60C35874A6219071FB7E491610176DBA20A3293B6BDC15FBFECA6ED9B97888077733E90075FC6C6DEB5F4EE326B8152046E39B3689C5C04AC4CE70138F7BD14A626FCF2637B49EBCDAB3002C27D9C96EDEFD548AC3EA77465921B514B84721EB8B75BDF027F31E9B6E5E20010B1A6B79E2285AB0675DBF1F60F61955500C1AFBB50C469252AC9739AEBBE78209D83C73760521D242D6F8D208109CBF2CCC5656E12ADA488DE17E03FB9D865F2FC72FFDB54621A663FB258F54D474D1AF93D6351A174A39D5F2BA98AC84CD68654DA67CE14C520301716D2B64B03A477A2A88C905ECACD544114907492318D1278A3F8F1CEEFC375CDB21C7EC8F4A1FF904BBC455F4F2A5DCC26ADD84AEDE22395ABAAFCF344C35EFDDBDF7918998AFEECEB52846522BE1390FC36823EB151AD2B250843E39EDAF2C011681D62BB4A02A8EC999C8B1D58ADFF9E9BDE47836065E94224529C23EB8677ED91BDC0ADB22CCA7E05AF174AEF5F879477CF1552D061DF28CB14E81470BE9BA0D77A7CE032675DB13117F54F9EA4671C671CE277375F580EAE03150FDE0B960AEEB5FF466BFEB15A464CB238707D2BE024B61016B98A66D6B0D8DEF3C193FDF35065BCCA948BC28723AC019E3618E77CF6E6A3DBFEE670AB7083D23E85D50647EAE84167FA22C6C8921F0D3A25D75A931754C8D7EBD8DB91DDA6ED5B54549630D6376580AC0ED1BFBE8FB4DA884E425DEF26832C05DC8F4078ED66CBD2855846E98578782539C9AA80DEA46B29448F3472CFE0ACAB8FC64EAF9ACA65A9529E62FADE1F0782B51DCFD33EABDC2B3EDB3353102E70F84325089CFB3D43099CD92CAACF9A0487E244A140E8FFC0885349ECEDC402728F493294E2A6F9C7665EA8C2FF343F651BC8F75582BDCA3AE807AF86C293A1B26FD850EA34B5CD7F37D75F0B13D7D837EA0C709F76625AE023674AA01621AEB569CCAAD76C29619C587DB7DD9DFD9222B7C5B871491B7F0AAFCD03964215FCFFB4ECF8B5FA8FFDA27DC9AAF56CFAAD270D8CB6132163926272A55769CBEF55F37324D84B24AFBF6DD8E9D4EB7DE1AFF726CF85A80960249D281D55B9FDD69C52B518E70CF1D3F69334CF8345F0CA8FC85F453068320B0C5A31CA1F1B32E43D6C3FC5B5FDB9FF4C6737C7B315CA5657473898AE2B32DC186B06910C3E4B3E5AE7E54DAC4811B860FD7073345A7612FB4DF86A599DCC12A9EC1DC7B61AFCBCEA6C122938B5944FB182266A4DECB83622CCBC08EB359A6D011E034097C34A8767BE6FEC9098DFA746D39FE40ADD20BD2CB59B00A2646B5A48B2B2086CEB23517621476E99D4FBBDCD6E6D468FE31FC326603BCB24C0B8AF2D09C18C56AD15B42A2FD72A90471D5880BFC16B1388541A3F18B582AF5D714D4BD7B5B73D7C7D9EC970CED3FD5EDBDBE2DB18960E0486D2B0FF08C43BEF34F8F3C4797C2300339945DF6F9A6B0')!
	cx := hex.decode('DE4E64C30CF4AA6C889FCD8B8C29D5C4DA1607B720FBFA7BDE4E1C5D5B733CAA55F4AF139B88C627D61EE5206786699E7F3400F576C0BF8E62004CD21C818A6EC03411F6C855F8DA0B7E78DF8A5C7B2A2038DEE5E2FDDF67EA78689463D1A54FFE6F7DE3B08AD75E1AE2F25528AA07CA94AFA4C2D089DD3E18C280A0B313BDFDD4A08A912710DAC4FAAE6FBF3BF72A6B191CA721CE7AEF8801A4F38B4FD20D89A22E4D521520E73BD0723CBF12DFE30C4ECF72')!
	sig := hex.decode('45F33C1F0DF0CFA587FEBE231394E160199EE47CA8819C82E21CCDEC53809A0DC3320B66D8F29FC294D87D0389AA6E25B375D245B20B16816F0739CD9FFE863A259CB9331AB93E3BFE70636955F352EDEA292B8CF25A8B865747B81FEA73B2F9C24937CBED62E479D654C3F1817F6EDBAE2B67EF845681A645A55B943F9A566616174E4698415127D5C8CB88D6D7311132E62D0F335B1F7226B787B0E4E45A9C2E4D93AB0C93F18FB0F0695DADF897D76187AEB2ED55A28A43BA7ED58CB0D64A09DCB70DDCAAD472B69B57949242A8569E4C732C716D07D341D634BEE84CFCF93C3EB100FF1CB6FF1F64BE283AAF4C4B842F0EFB24CA24DC244A70A7D8D9F231648B6BCA0E2E747A40E10F57D838048694033F24761FEB635BAE07C5E954D67D1EA5A243DDE59E1028E7FE125D1C29BA4F472F0788EA871CFEC58B854E487E8178BE8E0A22056E346F3CAF30BFAD0429E4E8B115ABAB3D7B8653BE2D12D0F7F41B2B2633410E3E995C3BA5437E4B883DC7B85FF4B1ADE28460FAB4D471FFF6B5EBE58670F405EA69B4D962D358C05950F67C70D661142020426DC32024E0A7CD379D08295944A5A7BE1B97C72A4849CBB916E2CF3B180E302F13EBACC829989DB86418B0D8BB2C897DB2006ED4B5D69C6DAC5E603937897F53D62666BDF30EF9231D6BFCBFD4C5AF57C77A7656D8B2E15A7B13E8277B8BE6DC16D744A465CB81A10CC766A8BE2CEFE5532213B3EA6EFD884214637ECABEB9F966699A69163A51F5661C6B830A0ADD66E3B931787D0366A4D473DBE69A4063C1B4EE8BC9E13CA1621ECD4EA78CA2168C96710BFD67D7D972714780899B71DD35AB693377C2521E73D6995A884E606E94407EA2B4B2ACD16C8C5FA7755224225E3C25CED4065FE5B1B5C343057A3793300C92F9A8F93F3E326C2E9BDE569E26749D5E601ADB3AAB673C3B5F54AE5AC0A8E67F30D0BC2EC144A20C45193D98F8F074FBF57986DDF71A1CA90166E9C3E07B64D280954CBEA0359BBA470DD7746F96B90990E51A47478EEB60210A44BEBA27C4AB27378143E029A55D8E83D24517D6882ED36ED833B85142B2F299CD1F8ACA9F0E144245FF409E9C09B32D1E6EECFDDF13F14FAC9E1D537C1C4B1063FEB0354DDA9D217687949EB933BF055D12BDFF4C9B9C162B805ECA8D63C868DB892248C4D1D844BC38939937CAECFE429904117D349F7414D24F7646D42FD47BE945F7EC6A3E6600C44D4339CA12DAF4D8B58A5437D90790C251A9DED082E7A39B305818991147598193C315D907CD7778D9EAA75875C2DA7F61ED5D1C2D5379A1BA7F23CA0165B2B3AD0C3D13FCF9C3B36C4863002FDF85884C3ECDC4BD9D39401162964C04ADA1B428B45866E2764655BF194E21C24607F120B56238A5479EE05DEB501BA09E714677C395AA5D1319D563EF981A753545ADA177E4B1A0F6A3B910E00EA6DBC636531EE88E068C229AB2AFDAD76DF51CF197DE702E081C786F18D9F28EEAD02B10D9DDF10967F8E64DEA3F51C4E72970E4FE28C361D893265FA22E573A4FE52154684191572E36000A758CFF2C459E23C9B9B1CA962DF4305E7C0789A2F00CF43A0F9E80A65D63B554F673BE96C6A36D671949BEA147A98AF4191BD8F61B4754039E8C7A3B3BDBF494368A556E49E1F0B4194E916B9D937579CC24C1ECD69FCA2ACCB0A8E63F13B1D6E1285402F72753672FC6A149D9FAE28FB7E90DBCEABD56993158F9ABDC2AD178D81296872CF444FAB021B1DBCDFC71AF3CE118ED7B4A8855D34E5EC5316C7EE7311327A28CBAF0B7190DA8C3C72DEB40D3DDF851D3E9240719074586A6FC0796882AD1EB5D1D7CCB3647F016CA91D7AEE1B6ACCC806D13F59A93D42CAB180682E4222E265CE90C09163CA03D6C63B2FBE8C53F542A6D8897E3D5C5B2EE781308668149CFAB81601498923B3356A1FC5E87ACD59205B3A789C488BEEBA5C4F2D1B70C8FC21154D4B6DC42CE16A93650F60F19D8D01593651BD60DAD6A1A3668E571344C3268F367A92521F383DE5F4A292A62C5031521FEE3E77C193CD8EFE5A4E69D5B7136E5E64A5C6EA6F53C3B3FEF95173282A673E54BAB8156CF459A6F92F75A3E14D62FCE2241172E25080E0225A6880967857BC058662EF1C7F9215080133151DCF7A897436606D53B2CD4904DA36A9146E833CD8F57847A7758498A6684EB4A99EAFC324B973268DD989E6DD73923A57D45A93FF16E2B7D92CA4EE484CAEC282A4B5CD59E0D559274327446376780BA0B4AD20024C0F1DB258A510D560294ED3A8504BDDAAC76A1BE72838BFC7D5779EB15D9A7D4E5CCF0057BB2124DB19EB737E7DD21F960B72CB3DC3FD90309C595A08E67D7B6207F067CD9D1EC23DF9B8EEE9DF2BA4E390DF6AC227926A73B78BFE02FCCE1E608AFE5DA2AF05C3A5BDD16966112724DFC32F6D32F6D39A026C8CEB56E347DAC45A3B1C0BECC0282F292A0B5ED2D36C706133D18AE2D252F8D9277C443134C78FF048167A3D1D94E0AA6C06B73EC7466CCC03528C9869B86A04EC51369EAA006BAE658FF49F597C72463EA8A8BEBE2BCD58C4D22951431B43C653C1EFFAEB01027FBC03A79FE7829F6B3B66A698D7396021BD92332EEA3D2DC485B1720B5BDB24341E75A676CD21BC650DC4D405D2557E874182BFE002A7EAC723565AA0FF2825019E93CDA672E13F26C6B1271C6A0F318BE29A9E1C2AD9893D2CECF135819D21C9A1C6A6C6568FB2C81EF15811DAB00718E8EB5C3C81C3E7842AA385068D12BFA5A952C84D00CC070DB07FFF3E5A9AEA57DA2D2FEDB95C1853216D4A17AC1F0C9D233B0B98397DE6264E90C96238EAB78FBEFA9699533B3B8B5AEDD59F1E603C3EE40F27FCAE578E982383D68C6936695B090A1545B1515D2DA5D66CA6FD80DDDBB73AB47C08771DF16E374755EAB703435CF049F4429BF7CC57698E5D674EB6423342B391C09903D4D82DCF52EF2CF339B5EBD8E948C69FB0E1CC71EED20E0F6F6A19E002F2DD727D0156FC3FFAAF9A8BD8D5BCC359A2144AEF4D7E78605891A7987FCDD59560F55E820E48405528D01215EC920273EDDEA684B01E383AD82FA3E139B3B946F5BC4AAEDBEE9755754D8C1909C4875F40EB846D9661D3857DE1DDBEE8DA72634915C286BC99654992511C8D756112D13001116E48ACAA952520415122D4D0232036AE605C73A262671E4AEE01B768E1B94D183BC5B06B64D3BF4B885CDFD13AA2299A853704F1C347F52B5ECAC30D97E6B0F4164EE9F4138F50BB03B31BE5E3535846AA4951B534265299A6CEA25C6F6017B1E50DA8360DBD347AFA0ABB2134E29C712750B74E7B232E8D7161658A78BFE2CA8CF08F55A90F90F8761DDEBE3CC78D07280F275BE9371678D5811798BDD7BF125C30675FEB868D7955B0229779EB83165FE5672A8F38100757105B337B7B2CD3D1D3201E71D0574D0EE8B219F92D1916BE2A4DC4347D0FD743B11153A00391E4411EB2B79FB5880F3B31A91B48C41FE1EF2C6F9D7B4D3B4E61C416C3656C50F422246AEF0253B917A34CF867FAD7D2FC8202D06EA7526B586B4E5B604A32F5B97170DA6A65103FA637A1B39F857414F7FDF9AF0CBF92FCB38DAEC89BE5D11328B9BD03E74827ED64289A56569A8F699DEB42D414A9F8DFA0CDC683D0A472F7CA0E84DD3D0E2473285EEBF55F696E7C26F88163CED91F5B2788563C04272DDF8F2409756461F4775E45FBEBC21AE145D22BACF71D630F53D41136FFB7DA0A55969859D3B76F87A214B2225A8DEBA0A9EABAB0C3FE895097A65F64F7661FD287CC52737D1A70E2D12150F2B79F42E9AC18B72F80BD0FBC5243F508F141F41A197FEEF24DF2644A82D66BBF4AB022756C33BD4F447081BC5D1416C138303E9D4D87AFF35E65CD76ACCD818229F99D169E2DB09FC9610066705CA25425BF7D3CA370709854B99E11B024F11A6560A3E0DD1E35E46EBA0A6F192F1D73F90697BCF8D9DC9735FF6FD5D492896121616653993ADD03CBA8E64FCA62CA61753E24FF35D210562E625DEBEAF7AA940E517FAA0CD51EBD9EEFC5DCF7F22B97F20F9570EBD34F35F3DB18A94DC11CB918F1B3B4BDDFBB78F50237427D7ED7309B2724D234E7EB632497C7C1939C05C0608087BC858744B0A1A837D62D057B6BAEE485C897143040BB5308D9077BDE0E8877A9B9B9892985FAA4A457DB8A320F42631516DCF746D3666683562629B76AB46500DC86E95785DFEA29962E6D21B39FA5E206C841575D8C79784C87519700C99D13812FAB43871CB0BD1A65242D0166D6313D87CCF8F268BCEB02D22CFFB683CE496499439C2DAA0705F612F0A7D61A8A04B41E528BC73E8A68F013B81E3E497327B7AA96D281D369D14758788D7A2B57567F3B95595C2960EE4597EC62F5F6F82DE7ACB34AFE2749AA6CFD4C26510F9DAA4750D4D95B37DA550AFA02D7D7ED8B522FE86C7212DCD55B7C45BC2387D4CA12F377FF01FBA6A5946A86FD192A7D88431409E6186F989E83C3429D1398586AF64826624988D48EB5D0F0990B5E0D1402C124C3CC5A84242B0FC487A13D197D8C5C560368B9729266CFF09C641FC9561B3F717DEDC8521F93936E08AD99203258E41DC9AB3C2339FBC919E0E0471AAD08DCB29FF6CAC5DE519D662307D21151D8796A3B0572D2BC9DAA8D565FE5B30649B2F66E5C6E18BBC7A0F48D507B5E93DDD9850BB6EF559CCDD40F7A8937166F75064253DA39E36916115B5618645E18C3973C5A5CD392963E393C803BE5845A06820EB8F8A1F9453BFFF7460F694EEEC9578E1808CC3BB7EB08E1F29D8261FEE147F5F7C94B65FDFE5F7FE2FEFB430BDF3A2417EEC2C406EAEAC70016FB860E505F5E44F67A3B5E14A395317AA256A84FC7609F570F3ACEFED41C934BF459B6FE5DDB39B5032FCE3715BA57C36CBB1968BB6C77C5369834BD9C3D5A9560595441E78831CC141AB7D80E290295230F1F4153B61E86430AEFE42EF6EABAB62188FB980269B72FD65929B5C4B893D11FB0F5F3D7CBEA475769DAB7AA9FA354B4E39C1FFEEA3A30E65A7B6997201266E90ECB5DC6819EDA816ADCA84EC739F0C188795E8A307636F848AAA715135C62D4CFC881358D34160E981F4EA7EF8C5A6D6254301863E86019EB4AC500259B5AD2DB169F322747DA3DA476FFC7C4E564E20710C111198A00ADA8D66C6947337C91F586402C73B9F1A147A98505CCF24823B9F7BA3BB55887682FB398616EBDF74C1D1A240D72624C43FE6A8E769D570AE5194CC59E60E3DB2416236187DD317F2DFC668EF4F23F9BE3831FED7B7A76345FDFB453B3631E236203A866508063C939FCACE9BC303F30A4C9BA76C12EB87921597CF53492686C233DC9EF45E293952A0836E1DAE197289F401AA581EC1AB52561A4F877B0BE1129BF1C9D088D4B1914C16276A6D9E618AD7414365A2719D0719F1EF8CCA60591DD23B18D9868F69324C485BDCC7393C2CDF2C634E29ED0A7192F7133990028333B7FCA8291EC220704027FBA21195F1FBC9640F4198B533A9793FAE53377B5307D6ED24EBAFBBC794059666692B08913018FA89422D6945FCF68383F4D2891E4085EBEFC8DE5B24A98664FA4425A1B62F2CCFF50CDFE81EEA6EA47636A41B82B292BC13997199FC088832545A23F7115737DCC903A07FC2BE52469C3C9512B46E42FEA096D4A485383E991860726A5AA11E91B8CC736D26378C74EE190C5186D030111332633DD4B9C630054B1289E887A683C45B775DB532A3B1C58741B80F4CAA232115B5BFE530DDA19C2FE84C19D5E31D7FF25D5F0A4472CF2AFFD02DDABFFF17782CDFCEA351C3847BDE52BD9CD4146D44CE623026950DB4E5B72F971DD8785D522290F938BAEEEFFC1CA6A6362A334EC95134AE0DDD7091271C8E0E00D6719484CBCF57536712D154DED7C6748C6217CA33CAC94D9C3BAD9FB13571DF8C3992A24E6063B9EDAEF439002414F710635B0BD261A7482ADD40CA74D3591DC12621B8BC706FF0492F80F60131A241739399D37D27CFCCBEE3ED13144EBFA5F832382669E81E3B68AB28C72279C859A1B8A1377828041DF4B8327C4DE1E0C9B3CFB648D2382712A8F011B564A806CDE1BA38F40A1CDE2D1C2E9BD5C409D76B25F77CC30A7D40AD645E8795984668E938EBA7E18934ECC20F4DAE563F33E76BFC1021A29A94371F57AD9336E967893DDCF293466255DAF00181BBAD785C6E081D8F3CD3CCF26E05EF7A9A9B367E48320B789F34334F5346ED6023F49D5CA008C2B8C866E09294F1880383CAE38EC563D690B34493544FBB80D5F7B361DEBF33D722D9D963015050F88F4554F7593A85F1E1AAC5C4FB4AEEE8DDDBC318F89DB31690434575ED8D6018BDCAC68BBB10610FA25B8E3CE7521911FC46D028323801F1A2ECB12BA7C3673F07769660CB4ED72A1B6801616A71C7321C06A0637F3D3A3DC3045A790446C53F4E1E85A3A93130D21C60BAE6B62F933784D10E0DB6D7772DBC0EB91CF0D7D90D0768F76709DEF4DC8577F9414A372EE8AE202BC886D8555486E8989B5C5F27B41F9E098CB829F73C97E33C22A431435595EC673EEA7EE6649828C48F2A78A063614227A4C4762AC1BA378235A785904319DF31FDC62C1A4D9CC60A14806F78ECA87442740EF365AECA36CB494541D4C39C5CEDE32690758E67561D8DD1B001BB1322CC0EFF5F45DBD62E8DAB75DA6EED8CB237F06F7FB3872DB6AD28EBD9245BA2E40C4328D88DE37910F4F8CF33CC176831D0972AC61726EC0766E3933A4171DAFEE475CF24FEEAF2C2F10874005428C03CEB1C8AD145133172DF53049A0BEF592AF8353814591BE9EA9CE693092F1CC6D99987EE4A9C688DA04E01B1BCA158341FACFD9EBF94AD5207A6EAB74B51500D8A2FF7DDC7B806994605F994FD1BCA410E4E67E8E3143A51D39A13C5F761587755A870DA14EFEC3C600747DAD49E7121BB7585EA9AE8E25A58150E8BB7288F349A4F637EE9DD6EDA296834192C8C4E5DA50756FB3C0F399B57F117171000831A7DD592883A31583760AFFAF907E25F51026E7EE89EA83C05A8C4DF9C1FBEA4C9FDE72E882E76C955B82E33CC78BFBDCDC3295F860D5BAA2BB454581B08447EE2AC774DFEC4042608C3100EE07BE69785931E4C6332918532421ED2B94D6410E9ACEA948F113FB221273E668E3163A1DD3DC1833F25088EEBAE3A280DB98AF0BD095557297897810B86B81297864385D4D0CD19765295B435018504BB387F58278A991C80DCB69F80CBD06D5D18CC440E569368A095359583A04A82ADA4665EC3EC7F5A8938F26D90BD8E6A29FAD8CABE532D011B9DA5ECEB4C9FEB6FF954893A00704CA8DD1B9B737B059685C31008C281EFC161DCD5279F90AA753F901970F41B5DCA7BD8CB90F1618BAD0B5813C76AB12ADFCCE91FFA59E5B6D37E2D39DBF4CE462DE4A4EB1A4CEBD239583F8BF2F6ADE1A37D47EEFA275837E9ADB7BC312D655DD628E857D6180A3E648661E479191CF6FCA305D643F3C1B62BEBDD8BB06271DB75D71B36D7EAE0DEA72549F1F26673FD566DE3CF80DAAFD90796D6C55E07DD22A08AC33F5B6C4222A2369B6D7A0D6F37F808DD5D4E2DE3CDD41E334F2D3F8C4D5853C19E4A2534C7EDD7F41ACC88DA0DC94513D6EE53209A2D53B10481563F49121F43758A470C44563A57B401830D2572EDA322655588713E92802DCF684A36EA7F4A0612A573618B3BBDDF23EDF345539761AD2FC779C2DC123F500D65E710F2331387D8F98118A5B67E92233CBBA0938572A01D17F8D524DDD99E62A92EABE67D1CE4B13BED634148A533C511302737E9D06E225B6468566A761D0952A2B22D1059C7D0A0F4C6113960D885290EC64C88F038A9445AE10ED0FAF804D69996690A70B1355361081C9C663F9315E7CF7127B8B0FDD013C9DA5DA61BBE565C870E6328B8025D8CF0C26693F5CE9105BA509934D3EA06F3C21738F68FA99E3282DED1B1CD9F5F24A98014A4DFEDD2B902AFA5003DCE3813C6640C6753E9F33B61297804403374AAEC9E0163A8DB2EC279DCB5C8A285A40B1FF66F2A62B4B8CD790F36CBD7B6854AC11D3C20E3CE2AAB8A36E04CD3DCED225B38F30486A8FDD79C40EF2583103AD20D3DCE0C4561D51A412AB5411C05F444E3A613F7CEB6806224987B5FCEAC4C0AB0043A22D5AB7C6F1020CE821FB302E0FF0F3F5F5DFDEE011822A313DDF94417E84030D74DB9696B7E192BC35E35E620D8A26359D1FDCEB91FD3096ED8D91B17C4854DD6459594B4161EFCC5804DA58B98E993828CE597BD6DCA010F70468054829923D15D0A1A2250BF58A3D062ED34768495E166B3FF18A59A01E25C623326C44963C17C79C425F9327C59F4249F44D3E2CFE084357883A0D7007DD188E4965E13C1CDA8C9EC77DC451B70DC91ADA52EA63DE58E7760524D149C643D9A828914EBF1B121302F243A9F3C5B2718A0986A4D2718B31E698FB329644A7C8D5FE1C009C678737650B2E314D4B64BBC4F90D4BDE0EF3E1799E554C908E074A6DE1CA5112091DBAA830420612CC518021A074DA4B78402CC052E07B6FDAD67289928F6718D31420AFD3D3FF83EE28539101990240C707277D82DD339CB00A4CD747C347F5FB71695AB6E79091C1C15A5D6FAF597C1EA09F3C4A55D23DE81FCC8ACDD4B2DF614722D18B9C5D89287E8E007301D3BB37ACC45F93D449124D2A0A75C920C58539852D5CAD778615FB6D106E159BC09E0769D8DF33DFF9CB85294C0CD847BBFB404AEF7F18159714F4AF9AE2D15DD30722EBC2D2B7494E9A022E2E15229DBFD06890F397ADEFAC18D5428EAAA31D0D1DF1A695BFF53D7BEF06EF8DE07F15ABDF4709A8096ACAB57663933134AF1E4ACACFF4CB98A3F61C8FEA26992C9950E6E10E03460351BAFCE660BB441E3419E32256B412E42831CCFE11F63A06AD39C66625C127AB08240D65EBE596ED20234B64463F6E0733BF945C9329C92E411D22F3BB07FE34CFD20023C74F21D9797DD9053064BE94206628130478385A7D4903A74CD1358FDE33A74807E76F27C3129691A6D9FD3CCBFBD5F1E3279964F6701D83E757F5865A14B020A62895F3FF8B2C57297333DDD5D74DCCE31960914828BE6B3ADD5D62430027932A2F35600801BE105F1984703E22BC961617B91AFAE08F815CC8B7F6AED9C55451DAB1D3BFCBBAD6D0A1C140F5348E971EE0EC8D27D09126662C3571D31D7612BBFBD8E33BD7467BB82969E6F79C9B23B3B827D94ED39CBD27600CB173A8C29A5B88AB661AC929F53060F2F5418B42DC50B9621F788497CE0C93E4856BEE0B9D152B55FCF9B434CD2E916D384835FCD3CFFCF08EFC4C54DA50B68089E5F23FDC00483A67C6D302F1AC45E162677F4EE2C233C49F08DC5B276E4F15ACAC032647FDAC14C1EEE18C4A95849F2F96038727D21E1258AF2D796022E10E8783533AB5D19C4BDE7200C3AF882BEE759B66E5F58A975EE63F62C5ECE3FF15BC8CEFC5D7E0B3DBF30939C0709AA7C48FBF2481597CB8BDFC0ED192E4471072A283E2D9397B6E44F23CB1BC9BA0F4FEB167D0F12A0EDC8B92E4D4069A448FD6E122FA7D6FDF2B1E139839EE31C788E80104C67DFD3CAB321EE561DFB5820DC41CC58502A400AB78E017D03CC129B97394D33B1D7FE2008D691F2ABD24D7CEE2EF9A244D3C8B6A9070BBB507545268C1B938AA48F8C0808ED520FCD761AE837A27262BD61DD5AF07D302FB6EDC5E8338589DB0E09C3B9ACF32DBE317B1007624C2C70505B0F42A8C780806BA276392D4B49ECE6DB836587FD208410F9B03525E6B431D8DB0C0D337E2EB8984AEE0A917AE35C690D6C24AA2465031BD1EF28963B2964A97B2E0813C880FF4A8E382DD4C0146609A195AA64DBBBAD81604D8B11FBC02468BD59A85EA91CAEAAAD4F6128F8CD0B458E11B0A2E2BAAE78A6B23E63C543EA1B0CB69CED38756EEC5BBE89392F4A9B26970C51EDDF23D9D32F434D876A0B2C7BA91456A21547CEBCFCBF056B90F48F01994311704664D197E60AA564DA81C5B8AD70EE289EBAACF37CD9AF9D23B872118E92ABF7D162ED1F5BB2348203DEA958D1180ABC6756B318844F0924B32203D0E0382AA1D81C749E4D6048CFCCF4EC259A9190D716AB29707A8B012C6C064B894D2FEFA5561C37BE19BF419BC88C82AFD53E649A6C6DE00B233CC9A31AE4A0F619F9E2C72B407781C75AD02BE182B0EAB2A7544245331368DB373DAEAAFC4F88FB3E2543AE681261F6E17E32F3DE7DB31543219F1D79E6EA49CBAFE608ABE0943C8114420781EC1F5F9E0B9C94FB08561B8376E7DE8846355DE74C1F3286FF7466B7F16463D10DE9654C424BBE8836732C150F810BA9A8BC110FDCFD959CCAFB23C6333A39CBCBCBA6FCAD5C9A67AA00F92E499F90279AA302F1A0D7E9643D3599CB4DF568CDBCB4FEFCD797984EFC9232D18F11F9A67D16B2F9E79E2B7F8A728F95593CB98A1AD73D62133FB028EC8C648F895EA9077385ACC647881D52EB00E14AC7D73D13AA4AA544C0AC9C901FD4B8C39A9E3B19BAF1F376E43ED5DDE8B681EDF7FA891A57BBA6B6E4610C48D3EFB549C801AD09F86E013B70EB7259CEEC573C219E828AEBA65661ACB5016B747F3865A6C51853C091B53D5485980EACC2920E6CAF918BA70168AC6C4FB0C6E1B84C79DED74B310CED201BBDE001DD23B581BD4EBCBD836D35F9CB43B97B56CC36211D9C11660B6BF35A76D35CCB2E3BAFB55DD56E608FACF26C4E79172B78BA9F41BDA3712929AB14D4546B258E1F2A83B7E7123D1BDFBF5305F7FA731ECA45D3542819B293EB9AA8509CFC0142E1E9A49A56DA58A155D8FF971160C8452B19CA1FBA59AE68754098B4D625535A61ADAE197C678E12F2A3955AAA6A28B06961AFA7F627F53E157C01265BEEDDAA1D0007E9898C0F1ED4EF7F87CBACCD4637D4C58B5A3367BB3E3F159F8B7BF7E6646DA93C5BB37986943C6E8900EE344DBF5F7066D7972BBCE7B80FD58425D0F05DA36AFBD3E551FA678686DF56FF9BA564A0FDBCFB72042B4A1C581946EB95BA020A8E6A55AB610838976BF3ED1BC477D20740D679E7EC62E390652900328F2DC75713ADBB01544B8AC68EF0E3F499E0820562FD67BDC9BDE1F8ABA63982BFC5712D71B0534BB525E4251E4FB907775688F360072352824491B9884BCA060651DC9C9BDC34BBA774815E4EB0117AD584E5DFBB74B837543199258DE5D3414724F99E7BE47C94B19E61E2578B01012C734F2BF2829A0ED375D0C1D74D74DE20147A0577F82E667DC42F7AA1AB794E94EBDFBCAF4D103C56774ACEFA383F75181BCD98DAF566C522814DAF6734125C8037E45F101847E8BA3C9668C45D8E82D4D2FF2140CCC0E1D26ABE7DD15C47CD98BF08FEB97D8AD3CEF63F0C4BF7493D16E3BF1485480B62B42BD8F7D51EC6A5B8C83036746D399F607CCAE7EDE14DC166CB22E53EEB3983B7154460722D4601C0E05C6D9264BF45A8390E37385B9CE1B2B565DD528EB693A932B24C9A0B464EAE56DA411E88E619236F7311AAB2D1B41C3D1CF8EA153FE134B6652A66A34DA0C456BABB313E8A287A2B4AFC4A8082F19CE4256ADD50DF4625969B5BFF89BDCB4334D577E03189A98EC8C87BFA1D53968AC9794E00A30CF25A7454F7DF3F99C683B910E28CDC0060CE7E12E429DBF70F8EA4DFF1152451068B37FBDEF14073DB7135A088949BA692139FF6A26FE0B5BA564422D47D869DCB18EE4353BDD719927D75880820A7FEF672532BFD69095340DAEE2E5FD8F899BCEC9EA320483361A0509BD1D4AC7F4C2DEE365CCF960EFD537FCDA4BC8D5B10EDFA72DDD56553249A89AFB590DC329D6A507BE8D863DB337702E66D214FCE4C965FE5E136B5BB375E37CE2787B5C71CE5EB65D539ADCCFB660A9D4232D690FDFE1C6D915B252DE10BE1D5121A10173F423F039E58E598B10F3FBC79300BCA7357E0741FBFEFEF149396B653D43DD12A8390608246C3C07EE45DF9207BDA8B1AFAC215BFE901324FD0FD942C3108B72084A93634315699B0DF845CF9311603CAB7D05F7CA3C68F576578E8A80505D93277B792F90D3EB5067764569520CFDDB6D2D3ACA895C922D9E329C40AF5EDBBEF7CF1C0AD0188F09E9B92BF081846B785738CEF4DF43363CAD744340E3959D1AA90467CC7A89FB8EC357C380201E00F41379BEF82B6CB27FAFA1197A8EFCEEA945BE41207305663C5E4454EF35EBD44259FB9C8367721FB78299CD418CBA9EC26D3CCB0879B376283A89C4170F03CE61690746FA292EA994C0E762B061425EACB8E990BB66D5EE004E5BE286562F121E4859AB3691145007200574EDC0D8571174A8D0DA378D386EA10C6297C6E0973B7250F4DA9F5316EA44C145DCC187630E8FD076BE140C88C05FBFC9F334959A64D47EA69A5E778A16EDB073CE540AAF7F389846AD0FDD96FF4146234D55C254FAADE2AA495B35CE5B2875086287F6E598D6015EDCCA90B923152BBFCF166AAE56FB69F3C0DC74C7128A971B63A8F0B2318649C601C4AFCCC44A7062962F656E836454E4030DCFC69EC81273102C59A3F1D222E99ED13D2BF61E577F29B73E8CA61A7C153E7E5A0F5E1E5C5A39A16268DE128277696D0011D9C9CB478973F88C282436E5B98F4B2D09BB08B070A51A9A645166F391B96E8FBE837B792BB8EF420A78601BDBEB048356D96789D9B18085279A05C93F35694DCEDD31438991ACB728116D86DB69A78DAADA2B6ADCE97D91A153528F563B9EB7901D94F10377B0BA6124E57180CDCA892BA7C2C0D09C0D7691E7DC4D17584A9C261BF1ABA05605A796CE038AAE23622D19678F523D79E17EC0113E39CF15BF27C0D94F6E5DD4F885D569943A39F50990825A793F6E0A57A9C50DF004DEB09758044EA51214E6383110BA62B6CC50C8C2AA024917B8C9F49F946F86016EC18AE171975477460531AC31735D7DF7614623E7DF77EE10EB34A14EDF2BB910A8B892C7C4FFF5DAD418A3294B305C9F7C6BC108479EE2828957D30E8AA2788998BF5350A89C23D97FAA62AF1A2B6A208E560965425C308ADFB1481897EB0C851D54E9D5E4245F6AB7FEDEC3ED08CE005AFA59FCBB47DABB4D8DFBFA8982CAE49147C2340F8405E4D521A3D6C55A6B2AAA22571E566DEF117432E650FDDC7C64830327BF1BB07E6BF64BE4BC5DB08547F2F5A55BF47B317EC09DD481F3580039E2830DB6AFC87EC7DF6F61277788AF1D11E08D4EDE85E2EB962F6721C73EC75F8FF1EE7C5A35831FC87627ED71B27FA98D07AC9A156E1CC3E188DC1CF943524AB466FC9345B65709D35F811C623D0CA469BD33E9F941279589E552AC3397933DD0D51D49EE115CDB472404D3D0D84FA1304B7048B02B61F664CE7524C81C16E89B624A25288A40508CDC9BB2B106E03346CD048F24417B8AC2153579F9FA1511B447B7BDDCC0E8A4AFD5CE21B08529BD7074649D6EA25C45D4833C2327083EC0D8D21A296F4622B5E16ED19D0E93131635D8E100DE05A213F309D4F67B68859ACB069BA507E438217C6E5A03D603DE8E9A737EA0CD985D014A8AB7CCA679935D708D5AFCEE19585C631D78514DD4F94374A56E6514D8720B08684E68154813425003F047CC97F419F680453F3DA090B21E8A0DB8B78343FD8375C1E44D27434232F0D38C1232DB10182D0FCAAFAC69D5C510599E3F7DDA99095B3BB3D71B96F274A88A889D2BE5671F377185C7B95B7E09955314BA9C52147595E289CC8D0D42D06D894E13A4077154A0DDA0EC4D5BB76C4AEF1676CD101B1873C36D9516E900273FA4768892A5E93E116D0A90251DED8805245EF3111D3C462E32C0FB9E329BED9D21CB8348962BCF8E72950DC84531056FA4D260328F4D7B1C11F5AAC696AD2D3D34135B3E3E2441791138A058AED7B094A981D020F4F246CB005F26F664896B4BE0C63C18FF1B9C53D102D45EB55A02F414C96DF7C6D5D866A19057C5A183F69987D26FD111DD0B6FFF3FC3CE46FC307FE40774CBA58982B2BB624FED8A64AC2693261537B9D379634317BE5ACF0A4A3977123DB9377A483C73C04E5654BEACD67E892808F51C30E75825B987B8E6852B741A9CBBED9642D208F7244D8214CB9E8F742FF4AE343885B3BFAB4D20B9C992FF0635F8B06498BD41A64326A4CE59493D5828F759E58E3A674C59F62E837F01F0FA6201355BA2A09B1851925A66D0264F251E01D1906ED6D146DB1C6516A88D941DC358031B0FAE9E7FB6D808032F67F4FD1390B2FAE2961EEC51932952A3C0FFEEB8ACD7E29950A76C2321175EF4AD8CAD7A3B69B6032AE21D94FA7552C635791D1D59AFE8DC4238061DB29453196EB8B7D794C80CDB7334D47FB8B66D2E21827FA4E04A24B7C81C42B62839594F4B5ED96D31ACB3FF16499E3A630B7446D461508A857E44FC0E90AA15FBF9BFF5743B88EF4E5174820C9CFD497B69375BF7F8BEEF4C089E3EBF0211B943FF6ED53D73022710320A5B06E6C264393F3917F70CBE848562501EDE7D8B3BCA14BB19E07A3480CD3264265C7001C3B1B7179180A377CB58730E79564F12F5D10182FC1EC632BDCED37C5EE67DE925D67430C28FA18ABFC2E7003215E4561A4FB3880D41BC5D7CA583D5C960402CE2F6B2518E2C103B53E2CFF94E804F6D47F72476256E2680CA685EF536BA7DBCD2013BA561EE261A8DA559765A7D57AABAC94E3D1FA1B1316A8F56EFDA81FD1657EA358762FE7F363D31BFD52BC74E730BD0A177115CF9625F2277E6242A38AD92554507CF402FECC017A7E9937407F25ED06C3A306D1D268825C169BE2ABD62291A260CE91125D42F443F96710A3F4CA55BECC0F74BEC44D80DD75B6E982B12660E6CC1C7FC3AE1156EF26D32079E68DE565141671571125FA6C00BD9B74B9B80309D2991463E794C8FCADA074DD0071E9BBD8A80DC953744012AAAB3E2D58EC0C3EB7FD46C5E052BF8A12E86E4F8347A7004C963F2DEE16FFBA71633F3554F1C2E3CBF71DD1F2584A38BD7E7D037FE73EDAF3DB5ABD292F93C0C1A816B99B133A2A7EE8E43409E917C8EA278DF7AFFB88840173E2A7DF81A06EAB17BC1853F42C96D0255B950A54CED71B3CD3153D159B0CDD1706DD4C4635C9F0C71ACA9C43BBA22BA977E4EE74B3630651E27EC8DE45B23A31BBEB23E6B762D9791EB185ABF2E4E908376EF38FF65E5EC811BA4AC45DDE55E9E39E79205C73332AE76161D0A0B785142D48FAA295E65E142A24760CDCBB4F5826948D32CC6C74AAE369B021289C5CCC2AE81933C8F22549620C7A513B07B0BC4CEDC52B502DACCC2C4280DBB04E37C13F4E005CF2659FB9957AE38BC2EB0A2A0E8FD25E1DC90BF582E1E08137FDC3A28AD8B3872FFBE55350C85549669AAE7F1A03A66FD2AB40C8F06911FC3B1F287BBE3E26A732F5B533F4F377EBAA2163ED895FBA49748A2AAFB3B1E5FA39B9E959E8F911A21E51FBBA87CFE01ADCF8440AB7BFF5AE73D625B8036DE0A159CA28BF4A0212016ED0629DE75C8F9568DE7B85CB5028EC0870E755F364C434EC34D165DA712AB6185B07DDBE1DAE99EA89C0589CB1673865906A4711584AD2BD9AF66B473AD6C41CECCE4FDDF222D8965C8996BEFAEA338D6E7CEC14617239060A6F9077BCA8C60726463F3BCB6DAB61FCC34B5A340E96F2256964B5EE5EF76E924B4615A4A370DBCBED2E016AB24D35582D7B4306DEF2718DF6C077C3AA45F53DD7A67FD8116207C63AB1D969F66C29CFE7C13F525F6B165954125985D0EE82A40BA8CE850E2111628D5744F4CB9362D98D94CFA942B32949EB0F55F7B3B27458F81C857DD7A66E933F409B575244185BAEDC29D3557F5E055D8F7E0F8D893480D276500A89FA20310032FF26CD6DD22DE2D87201CFE6E9D685A665654C4FD8B1ED49B2933F31404408264A2D3BA1DE73BB83853FCAD9D040ED18209F8DEC0E57842DAA3BD063D12DD1013044B8A4ECC0E6B0469820BF67986D461A7B3B905FEEBAE7EEE51AABEBEAFC4F51AD370FDE1D67F5130D46E25D9DEB2AD2A2CE2D51F73A4A7E50F051080C5AB319D741C7201C75AE181BBE457B49EBAB45D561A5C053EC9D21B5C8BADC424E15A116A8060042B32D1ECACA7EA477149BF4E2C7331BA90E80DD8CC2986FDDAA34DDCD8289D95912908151623E75709BBA7E7C8D69648D3A4B94081B243C06553B0C699882C85AB62B1D27170055FCE802FE9667D134FE262A72BC05B5FDCACC01C450D5B44CBED9BEFB7360FFD352D997B8AE146ACE36062A4DEF608A5BF735276A1C8B8F2252F533797C7E45ADC2653B8096C918C87EE8E0E3A1CDC9D9F3017EBA8CAB58B394A528F9F9B73F6158649A9A09E4BAF7EA2E289F50AFF86216EE954D672215A22D17F1F253EBBB00868AE0A3146E40A0E6FB8E59327B286DA5AE4F459CEE9C5B947A4176A8C5A3F64BCBADBD133F15A7BA3F62440DF8A67B785026199022D84CF01DA717E23C5418CDE5F7D4CEAAD03CE42A0B64803EB6900A10F4B3B107A28249E2413C24B0D494EB2EB043E0C827C025D27B022286ABFA9245D6895B6CC4095B7ECB4380ABC32EB71A649F14E047BCC6174FE7C323D1DF15B97B4DFA5A56265836EAE3AB06E2EC2591090E2AD3E577751B1500553FF6135EBAD6B986A09E61D5ABA190FB43AD5704755F1439FFB113FDAEEEC9128A4FFFFF22CCC650D52B174AC50BEE1AF046E534246E150AD71438072D8B456C12D6DC6DA13DEEECD94909675B7253A3199EA3AA453AFEE244DB1E98A922D126FCE6A86BE7314C08F4B3574D51EBC800257E7A0AA04EE5F99BD1E7977C3EC43FB2B4599A381851B76759592209940CD778CC5DD55E082F9EB8631DFD2FFC3DB3C2687A30BE6290978FB4EB94CCABBCF274E0BD28EF172334931D0CC9B815C2A6AE735900A3253BB70A148EC3188849159FAA084DB0089A1A40648AF318525EA46E3ED1BAD118B1D15B4F4F74EEF9058FF8C65C5FD3C55A9705A87A619160D4DAE9FED63DE72FB19B11B2E09FD431FBF47D53045BE16560532228EB14DEB065516B3518CE335647557F9D4A872FB2022BAEB5A0718E4FCA33D5DD7AD82049326FD0CD31A998F2A71A6460F646DF02E9C774FFC74EE12BFFF06D5A5DDF10A448749E20E4521D81FCB46CB7C93E54C350B8B74F58D640289DECA8C905048A6E5D71622018EB49A38F7BEB1735460BCCC3C0BF638DC91701A453625501889BBC13C897122AD03E3F2E2AD7814A8DC7ACFD8CC1B6C83D95CD626381DE3039A5A62DAD07E31F272D523CB9A6C6574FEDCE69E5164090FFF865AAB8BAAE934535B4B356D485B82031D00E75283CD09EB296BB4C4BD858B865DBC420800B960C1C64A3B8715AF030BD4423E6783F4B93B6E4E2D677DC809D146AF24BE579167B19D2A3C75855B36AD3B089E2B7182D328234321C5C12F56FEF2D7FED958E32D47C58969780AD887127FFEE9E42B82BF24A192F1B47E16CC82FA5E877BE8F75EA783DD871091C0045279E647C71956B63E1FB4CD13E9DAE0F5378A2304FCBCFD016A697004223CBA696F1C58B9BBDDEBAADC5D7C69790ADC9BA1F173C1BC8B2032266BCA019EB9F0B0884E68F3513410C53FFE1B790B4907AD1EA9AFD0E5DA923233170C96D01973C4D587644A30C60720CE7CC81A8DEF43702904C5907AECF788C4848CD6E52FAE9B1BE5966830F101AED158BE492F9CBAC6CD9F3BE400B7F4358CF9529B445FA2984A1580FA2EB8C22DE572B9D02F6B5584FDEC725A96B345DCE4693ADA9600B396CED6BC17ECB3C80DAA05AF669FE1FA5D8B9643E2210EFDD4C54EBF4A1AEF65D43EC2275F1752056A254FC28A3719F7A35EC77DEF17C687E8A0F684784CA44827B0397CF38CFBEA201CF0FC17D02193510D2F5DB3749F423EDB9CF2E7E15CF7F4C9602AF3F2B1E7D3A933E8AF1218B80510ABC4A21E348194C020149D59A0B90AB765BB4301C1B0600FA97A23A61C58F66F9A818477E9079056E7C72CE1921EBE807961FB5A11525CBB312DD701074493D10E40D5E7846555C377A21A2A92D6B94B7B6C7EF06CB7243BCDA35BD83921F8E8F54077DF68966C7DF0DC8DC510B910B1CE413E64EE5E8A7DCEAEF9D20B6F8D7E608D9FDFCF46F80AB3D96F3B901233B126E77C4F7D687029BBC7E1D9062AC6EE558173AF50F7B84D7D3D36CA808C8652C316DFDE021A51BE08A995445067EE51571D47B360622B5B5C3C7B7FE9E254B587D5375CEDA31EE8FD1A496F60002AE444C729D2E8BD286B62A7D0BC43E91BE5713B88C9512721953C61E1DA0B87D469DAAD2AF7E6AE21C2391E150D5DA364AD3EA46ABFD34CB24F2E2B91B8E94FAF99C0F20C1DF6FD81FF028B6D04FBE0EED84CD7F8CED0984112A884810495C11548AEB859608AE90553112CDFA0CFECEFC7B392272694E206D0BB078AA554A1B1C9327C30E6256EA377F2869E775BF131B2D8F50CE60522FB0942D532892AFB078BC1CCC3C6607DF37A1DBFCE78E92ADE275986630583870A9EEB86B658AC371FF39EA83C25F510E52DE5ED5D0C031481AF13DCD2F3BD15BD29D5084F65C175C050A7647560F6169A489469B047FD370ACBB6BFF34C896BBAF82B5F032EBF5EBEEB4E25F4EE704967081A43510B186E35693593D5B0904F51FF885FB3FC5940523A64CD0BDAAFE13C6DEB26F1C539BF15A672B56961E41195464FFBE7B898E4A0B0818D33319994BBE972A792F8C208742AB042E2452182862CDF7578EA78D52ABA0BAAD79774F51E6F7265CD5C38CA2926CAC62BDC6FF1741F2E36FE552645CB3683F9A7D2DC12BFD8A15F9346B3047B2E14B513A6D1934013338200425E947F8011323C559072FD9EB838E263BA075B1D207AECF29B53BB5A490F7A31C5992E21856771654EAE0705D9FCECD866C384001ADE166EFB028190F087D17C29AA87D1EC14A3ADEB40B1B076548502B9DD942405D93C01FDCE562AC6DE673EB6798F333CBB8B110A0579BFE0B93AB6B927813E054C785393FBF10E32D557C26697F50EEB850E0BC52FF977494B21554782BD96D341C469AA9ADF9258A74C6E0C0A0F9E71BC09532848426CCE1682342D7C8CB3F4D509ABC7B145E6CD51FEB0F06A0F2AFD53173CADB5D11EB44187A59ACBCBAC953766758D99977996FF685C0E5F69A4AA3333CF9AB7D97C62A6869B4E6BBE6C7D204B78392DC8BCE9ADD8ADB3AC6B0752E153043427B44D154E5E2C879A38F1ED0CC2A500203B976EF303D8A432235BEC8E117943FB882D90FC346B1658E954767772C68FA55B58A7B463BD6281543A7E7444F0FDD4140D5FD8C78A1EA9C99F27762D108ED4EFE91E4DD269D9AF01138BFF6EA6AECBB80FE23287E2AA3E6298867ED88283748E21DB6E3C123662649E124023CF6CF7902BDB03935FC496BCC5B4E5948BA167BD7C2589CEC444D37594EE9E05F032AFCF2205F2F1B6DC2126F2AE499292FB8F97E4C61ADAFF16904296BA78F584CE30210663C25C83475F399899F0DCEC73FE7CCD3F2D5656018ECC491CD5DFB0619029EC8CFF95A13C38AC7172135E0034DB24D59FB6EF57612ADAE2C66C0F634E500EE5C1938E987C57E8D124742A333F48EBED00596229805AEAE38480451F3827E3DE1FFA5E6B562FFCBCEAB6B6666502851C9D162787B235687433A567434D61DD1921A0C5FC6B46A9728FF850B74C856A3046BA5E4050ED893DD7B5E7C8EA9A5DC2344D2D3BFE93419C2A3F6D1E761C3F3E9E0EFE16838694D57EC3D5F9027542163C69A537C8A92D602D21CCA1246C0D03B1E549551C93D70DF28C4240A180023179CA7137F4F4403EF7F0692804D78F68BCF3C536E781F4281E3AC276A06747A0004E2F3CEA8F79D5DB17DEE0BC632C95F39B7374C988398EAC6D7F648F2CCCDDCFBF9C2D46A520645C6D60A775C3B423C8AA6CF367A4E0578A3D91D1AE8A13A9C69B960437DB8114E125478068F37BCEF4AC48FB5A06CB5715ADD19C6F3C4EB90998A77E492F1D56202CEAABA96A5D9CD6AC06A1A4535E294EF4BFC3C1116C3FA16496DF058F841C9D87A04F79EB6E25467584F5B1E002BF31BB2FE2F407701E2EC7483F0E23B788ECB6E48FAA1E6B49A729D56375D0DF8926334308C547386C6290C2768AF0A8AAA5D3689917A9A59BE4517F7B988E670ED5F85266F82FF76E3506814532D8F867008714A038CE776F7E2B8C9A4C148C7E8E7BC4CC45FDA27A0A5BC114FCF88832B28C044A41D70327532858976739D8283F2D7D7ADF706D7777B57AC5A12574F34380898B85F1112CD5530FF0DD3A6CFE130E0B184F91AD20F605AB41CEA344811E5606BBD787A2BD323CDB70AC408DC7A3D92A429A4CBE879065AC01D773F7B678193D21E5B4049977148594C8A909FC8E272F1281DD24386C518E694E9D1BA3297D7A2C07249275D743B46512DB3A12602BF5DB3CD7C8F113BF7590EC234801823FB62658E092D3050997370BBE057EA30FA50C075F6A5D8A6337D5E4D3B7DAA516C37CC166A150F98C089BB7D54527CD19C9D18459895EDE82725B1D65862B1E3363A0D9A3DA7DE740EF0E699EEE6180A709286C268E8EC6D80412F7EBD53A50B92959D43571AE562069C908DCCFAA491CB5162E553CC2E9EBF46C6124E9EA254A71F1A5E168712906D7AB550BF2B6CB6D60E04C8F2392A0CC9BB980212DB515CDF7100E457C0E4DD3AC8FC939E5E3A426FB88AFE7334007A401C835BC96E838264D0BA8AACA783CDF8767B74C99EE590C3CBD0AA605FBCE8EB93E9F5BB9B184D9EE8C6E5E0BF8C00D39EA6CB9D8984D6B01669218BC62347FB9B15C9970B847C9A08008EC3FC329C7282E67C44ED844856AA8A8A80B2E7D81C9AE6607C3F61EBCE95A5438470AFE70D609053C5BB0D4D65934A73600F248D4C2BD56D4F5DC6AAF00580F9DBCEFB2BCDD7C11098148FC5EA829AF38F480424E57542C376DD49D6813E1F0740BA90AEFAEF590C855EB878B505B70025089896C4D251DCF7464F187CF8C0A3D6EF605D8888E7947C4038856C576322B2BA1CF3E90035B88EAE2469FEA2D36456FD1FAE1ECD89932080EC50CCC6062EBC9328041FD8C08F235CC5DD24EBF237947D46E0C6E34BBAD76F71C748053600D08871AC266667A46DC4AB10741A9CB92846584200E497A51A59E03E06CFF5BA68DEF19A05C954AA807DB4C82E4F6BA8FCFE59F1252740828E030DA9E441511F2A78B13D3619AC9AEEFEFA20257F59FF0DFA06005645F0B7FF1C9FBBC99F39A13A3755841A7CF70F39CFC0087954C1A7ED0E36388628038DAE4C2D256EC7E84FA4A32061AA1CD04AF0DD003E99A0FDA1DDE3055C2192CB052E92CB9BBB13808A405CB50D1BFEBE3EE1FA38F9E91889FF2B82DD3CD2D2CF2F374A414C26A20F72A4805A9590977043F854A876518168AF69F43B2A01BF870739D23B9EEF5720F551C0AF918BE9B22A400E7E720660BE200B50ABF2FDC4EB57BD7C3A3067C0B744389469C571DF9D330B512263FD589B55BFFD44D1C407EAB6301CBB59986B0EA80FB146CB9FC7979E1CE8C86826DF3FBE314EA1250C6469AE84C55E1A9EC15AADCBEA4CE0AEB40CE6D2010D720B2F74B34C7DDF1115386635871DE19E60E1DE3B8FC43DC709970407454606066FF7064C07334C74A479484AD30476C64E6BBA91F8D9291FD198E9B2FB0C6A05C86F958F534CCFCE48EFEFEB56D0608D82462030A024B9D43A5919FE068B054E4FBC7A90DE9136A1F498C2F572ABB4A91665A971D527F19F11E4ACA0EBC72E03735DFA728C08D5D1BBDD53A0FAEC3A947F39FCBC4CE0BCED31CFD6E5DE960F10EC621B1CAD93F78B9A305A82F678EF4C2D5A6BC4D2D62C58066BCD3811235F1521397E9DD835E0C7D878E1FF96935B3FBB48ACD0283D47BDBB6CAB266EE23FFB1A81E7112C3F5E4E692F133FAF1531CE03E3C9AFB6BFE89B2824E7B3CA515D0FA9D4A74B354CFBD0AAE9BF3635D0A23441DB1F32A77DB4630134B7A81A6E33568DAE70F85701E5A920FFEF927463E16B60C58A211C82D1DDD448B0CF0F86553A37BB4A3F059A9F81492712260E37DE4D3678B58416B3EC07C364B1CF8BC3A033CB23235CAEBBA135278DF1FC368ED1E80EA6F017BE64FFD64CB265B70033A08F94DBDAAA700FDEB669E1FC1C6ACF93F7DEE2B0B31A43AD6DE01753A631593DBB2BAFEE41B9D5D318CC250DC5DEEB48EE4998C2C2320C2D3D8CA6E32F0F68112F42CFE1EC467DD7D90A0FF6E03008C628FFBA75B172454F35E63EC3ED5BE230A40E51740A85C91CDD0ABD44EEB057EBF08875B9590DA6081A70F1CEA241CFD24EE5B388F09FED5549B2FFE73D2E02C2E9DF0B1AB07A39424731F06539F7B210CB0889306A03B34ADAF4E84CBF22A0387802049EC2BCFC95514A560AF53781DB9061282BA662DA73895CE766AA190B6520D06720D8FC0FA8BF5A741194ADD6DF957C8C30D29E575B9FE5EE6EB024704F06CC4F1B2FDDD053B4F4464ACF6356E2C6E4EA41ABC4A12F7BC71AD362AF657D22EBCDB363C31B1773E5B8562BAF7CA187830F1B1AA20597FB8D8A0DC0CC6428CB577AAE8E9C17170283EA2689607B6AC6AC2661AF2580B21574C89B06947EFCCF4DB8870E5C3EB7ECC5FFD86B0B51E72F18610D32CB14831E9D787F7491B7AE593F4AD6F9B4181B2D2CD3CDA5C82B1FDD5594568D3197275975139902F5A5720643BCA23F542043735CC840BF5EACEC5C1189514DE081ECE6F06DE4D20042933395B3B45707514FA39C5009C78E28143C9F997E013BFC1DCF8E55F0B399EA4A62288852F33FC8C317DD864811E2B3D237719A5B8C33F6FDF00B06905F23D2F4E8836825F5ED81B0F69A366CDC5463889B391BDF67176E63870DF39C3C9DC2B0343BF69A2ECA2893A19F569FED8DD8FF264A10BB0426A6851B42D4668DFACCF60D2A7758A759D2E6813AE47CD91B2DE4053B2EA372C2E94303CD753563373FBAF747AC3E8A5068231C8CD227B811C3AA3A63D26FDE2A85D9A27908E18E9BC5AD961018F6363264C4B5AE4B846BB14629984CD78CB0C298072887271E5A81244C779D8725824BB8D3AC99B4586BC17BBE82F1E16689A860352E545A3816D1B2CDF22300D2C428ED618F6107E8395A2BFB44C8BA75ACEBF7F2718B84020EBB86945D465E7EDC610598693E44E00C0F11655675052FA1596C912E84A0D15018CA5E561EF58E2B6C48D7BADFD9D36A85A74E27E30E4DC7FA61DD5269E64C9215584915A0C599A7F211D7088BB7A00AD147C4E1AC9B0FDF4762E4623AFDF9037EADC3CA2405D82668F2E03C56DAE28447A66F94F7AD44333652673A8E55F2C167D998C1B921C6257ECD99D606622D1A6B7B06F1F2E7066FD2772D4C33DDC5C1A5FD9C1B960B58AC4A17E4BA79AAC58B8CA6966DAAF14D61B9B2E77E6610A0E4230E158483A04A851E8F1F63EAD0B8C26E3982F0598614BF1F202DD41B0DE21E44BC562E203031D71CBB7FC00A799F1B1C0AABEECFABA878F010EF5F34B964957BA18B52B0A5DE99804B52CED098603F655F3F4E383A631605F5D8987FCCD2D601D5879619B0CA49B55B4AFDF195574068C40A71D5B0215AF8ADBFEA03FA7976AF81BD7D5487E84789EA0A1B41A55C2E26611875D260BE02F4AF2E7A66D5312C9E561B6CB213BDCEED28AD7EA890C213DD92758CCA36836A77D5F1017C1AEFE1BC8DADC12D5ED64A7815A56F6A355CF9DD25B6DE370D4C9EA86F97913319B0FDF729729EF7C8693A69C6AC17C3EC8ADE0E530AC9F9733AC4CB6171239E113C8D7C7FADA46EBF87B203EF412919ECD5C03439A16255613AC3CC1A829990FCDC1369CEFE6A5C9BCD25F7B476364B9A969813B57E1CD1069F3CA4E959A7BF1718DCE971084ECC6B7A5C2889053F7EEBD990889BA1E15E6DE7A021140FFB264C4D32AB34F6CCA93C0103487438FE26313E5FC3A333D754F33F33BA588320AC7A4F3181CA2CF234E1B8A5B831E9AB5DAB35BC7B826E152F300481DB7FA74BB795188517B9B5EA86A91E5E9AAEE6C0B8E1A77A01506616B5A40CE7C67F88B5542F0EBA5E9D9E4365AAACB1CBEAD207A93A9CD339924FAD5E464969C0CB4C06D9B8DD9508CE44BDC8A4DDB2A7F9B30F5F6122D7B106DE342C3388154CA41CA612E77B59531C1112FD0999F641D6E165490B692F')!

	ctx := new_context_from_name('SLH-DSA-SHA2-128f')!
	sk := slh_keygen_from_bytes(ctx, skb)!

	// signing with custom random
	msgout := encode_msg_purehash(cx, msg)
	outsig := slh_sign_internal(msgout, sk, addrnd)!.bytes()

	assert outsig == sig

	// Testing with SigningKey.sign API
	opt := Options{
		// non-deterministic options
		deterministic: false
		// pureHash generation, default. can be ommited
		msg_encoding: true
		// use testing entropy, for testing should be true
		testing: true
		// set the entropy to randomness value
		entropy: addrnd
	}

	sig2 := sk.sign(msg, cx, opt)!
	assert sig2 == sig
}

struct SiggenGroupItem {
	tgid               int
	testtype           string
	parameterset       string
	deterministic      bool
	signatureinterface string
	prehash            string
	tests              []SiggenCaseItem
}

struct SiggenCaseItem {
	tcid      int
	deferred  bool
	sk        string
	pk        string
	message   string
	context   string
	hashalg   string
	signature string
}

fn test_public_purehash_deterministic_siggen() ! {
	c := new_context_from_name(siggen_item.parameterset)!
	for t in siggen_item.tests {
		skb := hex.decode(t.sk)!
		pkb := hex.decode(t.pk)!
		msg := hex.decode(t.message)!
		cx := hex.decode(t.context)!
		expected_sig := hex.decode(t.signature)!

		sk := slh_keygen_from_bytes(c, skb)!
		pk := new_pubkey(c, pkb)!
		assert sk.pubkey().equal(pk)

		// sign in deterministic way
		msgout := encode_msg_purehash(cx, msg)
		sig := slh_sign_internal(msgout, sk, sk.pkseed)!.bytes()

		assert sig == expected_sig
	}
}

const siggen_item = SiggenGroupItem{
	tgid:               1
	testtype:           'AFT'
	parameterset:       'SLH-DSA-SHA2-128f'
	deterministic:      true
	signatureinterface: 'external'
	prehash:            'pure'
	tests:              [
		SiggenCaseItem{
			tcid:      1
			deferred:  false
			sk:        '3BF9B2D4368C24C95278BAAEDA5268CC38CA32BE3DFAF435E9400F18EB3ECF812AACBC8669722400423D9CBFC5E3FB9ED5717C0C9F35FB62DB7437F5C5D4D387'
			pk:        '2AACBC8669722400423D9CBFC5E3FB9ED5717C0C9F35FB62DB7437F5C5D4D387'
			message:   'CD620CF74127F8240E9BED33E9348183C2C9955E8383583C3CE3934B53A6F30502DA5CFBB89D58360C0C9C40F5135919B004809DC4720E2A5EC495995D0430AADBE347424E328743665AD092ADB601D17DF14F8351CFE8491DAA2D40E1BF90DC9E49F7F7E5D70A0088D26CADBB2CD58B057659EEE0CFF4D3DA2C1A59321015D3078CBF82420648D6DF305345A2C37537036050F79397685ECC3AFD2DAEEA30DB170F703164D8EC556DEC86492DC00DD759C84363EB2DE277BD235B2F5BB5C366798006AF9BCFFF47C33C24750F2681276959E37150AA5C1DBE0C016420B0919262966FAFE876313C39940D474BA083BE887CDFED4725FCE830EE25CC0C39DCD1846F1693E409A449472A974C928C0CE4D80D9DFD811502782954B98CBF7867D0E1A0D457845CCC25796103499E253CE97BE545740ABE7158C79BF0B02F1EAB4A743672CF7587C91D82A8BBF36DC9141A05E9AA6BC3DC06547049DF4E7A4ECE35557113B34042D2265008511112E1A1A7EA6BFFFE5300BC88E9B21148AD1A26D3B9CED50F71FE8504E7FE6B8065F00782918D69A02187042B8184B1C546B924BC88B6011A633334530C2185582C3E0D9B785802D2D7AF89BAE83943A55191256C5797BE728B7FDA935F404FAB42ED64C42A03566C267C5446298C993EC794935CCCC7469002389ECEC4284E2CF5B24782780A3AE5EDF2349D28C0AB294E9EBCAE6C455E8970DCCE65E8435E5B197D07D4B6E8DD8443FFA22A50B66DD19E8712228368A9FD86FD6A558E7EE48F1D8553969249B161C140171543E587DA325DE3CDD37BE06D14991D67499EC45A15E510D8909F2E8155E69E64D5BD97A465B3F453D8FA752D5DE436C0CA064760A5EDD3DB89EC8E26B0BCC848A83D514A5AE86E90FF6947E9C199C41FC5DE3E1D2E47A22708F28CD344F3BC20E436C72204FC9E092375A74714DBCD15C0D3196CDDAC7E6F605546F9F19206A6B15CC58FAF85F2DF4B1BC9ADB7027C4EEB7E654A996E7CA9C576A7F6DBEA25ED225F49912AB994261DB3DB5A5544E6074C22E3177F2905FBEDEF4843AC109226761FF19E0AC971CE95E5739F696A980DBA54076E109B0C14FD535A9C87290C915244C4EE51A05B5490F3B28B3D024F488CCF6DB8A2E56B3A0D433E651D02C24771B1A2B8B224DD270CAA537BD619573BB9789E4A717D43F5FD76132EC868FEE46F88A5943E09C02A19DE35E5DB69B1207107CE1CE632D01746E1C1724FF606428F2EE4873AC9438894847C429489D6BFE96225CEAA8E135410E05E829155AE9620CA6EB2289B8397D679AAF986E1F7A46353C8FD8C260CFEE00D23BE6119013F7E03238C2D3A12B260B2F5B78DF362349FBF9B92942C9944569CEC3B4DE34ACB3137EDE9159763FFE65C2A266B639BCD4971A2ABE532766BEC39239139F80F8AD8601B28C1ABA5416A80C50B98857D7A2E26345D6E232C4C60AE94BBD8CE7FAB68C2ACE8DDCAF37DCE10CE117FD71A81F4FB60B9A4774D8549F9F3B4297351399244E2B20771758FDFD9D4BBA875455363BE2E2A0812F04B74B359535AD256A3CC7787C42A7D3F232668CB94C2C138A34C4D877F161EB019090D2F47949CF8AA6D977DE01992A0EA3D4548B82BF958A4FAEEEF527DC43A4957A057CB687D686E21F78E1B6633913C9F0444516808BA60D998C4FD0B19A1FCB3E414AACF40EF8297B0C1E65A313DBFEBFA6C1FC0ED2E6C4B260C58FF001FE2DDE84DA3F37D370B24053F96740586E5F0C4FE2AFC7FE500880727064C1387D74736ECE1162D84E925699EA5EEB674722C586B87D76718CACA64D177665C75C2AB2E4DE978B33D5C4BD5911549AF645A7F8E63C1D63205941F6494548AD0BFB77EE8555310F3018F1942B9DDFB382F5FB85C482614F3AB00815DDC7943579F05B28D4D780E1DB6C7B477B5823286F2FBDED8AB29D57244CC616370C7BBB507CFC5EC63ED340D3764861D9858C00D64F225982F4B2664F1167B828646813CE54DD0758F967817940E23D18EC689BF4EE7AAF203A003D8445483DC05C81B5B3614E421180FF40EE4293832236BB874F3804AA2A1B750C96FE98584A55D40CC40463D473B7C40988A4BAA546A72C1CAD8283946945CA1735B1F9E59A87E598E7DA3A5E435919C2CC7DFFE432BACE90D432D03FFECBE70E62B72D9D7A90878888ED500548004F7DC2725050543CDE534F747612007E8647EF725E92C6EC352CCE4421010E0E054A44E0BE7503D670C159F479BFCD45CCB9FE6E134D5A945E70E76426C4FE2847B9243367CD3874A602CFA937255D2C90F5091F3955C7398DBCADE6E9B9D9306A8119C6EC5E3AD5C927B3DA76D8410C57D12E000558A961800081A2A2F1AC69ED36717831B50DBEF51E77E2C7473A1F5F40D89613C676EBF95B8BEA1D3FE4311A8B21B0E7905D306741C67C44A2CD0BEAAED28722B6E50EF769188EE564F0BB9ABC85845324BE21D80B4D08C57E5511EA714F0DEB7EED900F74E595C2253BB44A9BFA99C4A77D39ACBE061056E483ECFEDAB421294B4785464A2BC06E6ADFDE1B93FD495B43FCAE926849330433EA2B4553F0A203475837E555EDB1461FA1F5F10A44411FC930FF8CC77871833CDB340B61D00060D0D86FE51D129C4379660AE9DC6FDF77F59D15645172EBB73D54F7E2313AAC1A8BD260E9CC36BCDE9550FFA32FAED824CD65361DFA9C3331B22C1BD9F131A479193A98A494ACDD3BBB1FF084B4ADD3492EE923D5A3B5551476F586996277EE95E5A44102F8070DF14AE9D34FB0AA2748C58E41DFC78A2D5A3D80BB929E18158E5FB13EDBE698C770C8FB6FC11F92A5228824B188064E472480379BCF77C6ECAAAAF2E255DCBF6D7706482E1EBEBD81D95023698AC2C08142171B9B541FDDC8F71A1E7EA17BF555F1AF844887806E302B8BBB9D30CDF6C929945E5B32A11CFB4EDFBE8CEED91D94ED6427718BFA1590624E4C710B1C98B5970D57CF00E2CA29211032AD20C08E67FCC6B9D9739DD671535F3DFCDA4E0B817CEF4D7D411A5BA73DAB1F526B78EF904B16BF169E0594E48A98D95C8A07C43072AE160060C98EABDD57DF0872511A2CABB7F49E7E7E2F82EFBE46CFB628FF1CA381B385A58B583FA53D94CD987492C1588F85791467C22623CB9BB90923D97215678D051262BC213118F630A4434E8B675FF39FAB04842086C5F861BC8958AB7E3910E7000A114C2F208DA89848EC1C2D484261DF57AB265E8D0F23BEEB41BEB19E89806F7BC3B9B1C2E7463AD2BD95F9A74D0E480A49F7C97052D3B3C31F1676B87B45EEE5C37A568A6C195F74A6A150C2F6DE01C8773CD4787632E62A341DEC36CAD1840E58F0755EC6BF371E704FA348FDE7E10B5D319A0F5437D648C91D39A337CFB459FA4EAAD7D96EFA013C38B05C7BBF377DC124067F2B7E5D03D85EBDC0B06357209C2EF83555A22F53A0C57DA14BBE9776EDFA168EE04078F2740089F8B2AAC6A9D9FC0B03362567D7A2E6CFA460C1145247707B871D211CA7223E5ACD89D24A7069EE625000EEF7598123BFFCF79B20CECE13CAFD2B20984C4C1BE22D8EE90B62E3B73F919FD276127D96B7A56D68B3146BD9A685352E37A980023276F164F038D92D55BABF8CA874A9002B52DA184E8E92E3827F21E4803961FF2E38571F1298E981CDBBE755F7EE58D869B5679998AE4A998603FDE9CAA6E94D00A77AF15D02B582EC62C6991828E78058EC8B698662969939A421D81BD5E48454FF7EEF7EB1C4F52EEE0C2F47843DB7EC09BFBF2B3E3C7F86E9A31207E460F8820E1D55D0D39A18ABB697B2E22D82ECC629BC8CDE769262454FB308CA60ABC6A0EE5CCA6103D198869E35BD9081BF49E27D82A3AB01D6EED87E59A27C20A6D17438449177756A48CD678EB5656AE0AEF22F2971421FFEE58FC43FCB4C9F0015439B288120A1691BFEC4B3A9E766A31849A6417C35FA7C9CB96542D081591D8101761C08733A45339B6F7BBEACB84AD2A4C1245A10018B5FA39BBB65E5047B6A836052223957D97E00618DC14A102864CB37E50CC390E153A845604CA845951920B5DEC52D160A89DDF7FB0165239503E863BB7A2DAC2052257F4833E1B775FB62E2F4EF2400D876A202B8E3F316D2E08942041E40F80C2594F2D5F59CBC9C96EBFE1848142E45EC81FC7229D1C5550B64D4E08E4E51E97B2B090D79FD5A73243C8AA9581247B569C042703A73373EA27CC3400FD0D91195462A8FC998163EF226E5510067C1DEB4D4C1575FE73FA5BAD295802C4CAA099D8B1119E0FC9A3B17A2676A18E20147FCFF9CA9EA76ACA6601B7C63C33DD15990FE4301AFCECE418EABCE0C9D9FB1273658BE0D963B07D09CC0E8AF3E18D6E5BEF4F9DA1947A0BAFD32D4E257497748CABA8C9A13904E8AC85C595079BB74639E154604D87BE1C2F2D19DE4B5D03CF611526AB27C650AF509D255FB0A938C9B179AC2843F88AB256D08FF2E85586D2E4763E406469BFE50A9759D73A14ECBF1F0234D22FE745A0558B14E7AB5A47A9755F749C6858CBE64BDC108898E03E6BB73B4C30FFFB315812A798304F0BC11A20F2B7797FA4FA6C3333CD61405747EEBC64F36D74689C2CD9F34063C5FE19183D50E0E0CEFACFABA8C1989B270A4C530B5E2F6924FF6A00D386734F4FA32ECCCEF56C8CAB534DEBCD176CDF696FB34C428F07F3CAE80DA9DD8B341BE69CC215A1020ADB578FE31251FA5232A9488C07A259EC11B8CFCED9D0C31C8E669EE520491527F67655A62EA1BFC399C1DE6DF91A9ABACBBD0C2AC9F88031FEBE84D2149314101742A7A15D25A91DE398C65901C1DA1338B37934592C6A9D17B3CCD7BFA35B5F1BDF2FD42ED36E44F16657339598E4CA96447670F22FEF4616D574CC6A9A843BCB5BF2E68C7057AF246B63497380728C7F367243DE27BB0DC5BB45868293B055AFCAB30825640008875597AE3DB5025B5BF65F1BEF33067F63174A8C79DF04BC1AA1FF76DCCD83DF516177E4A61F250F48BE65864FCAF6AE4190D6A9435269FF393ECD62C54B1AC17DAFE6E5E247103AC08DDFE3DF3DFBE704C4C1F68F008E38475A2CB759E69D28A145C44BB2FA73038765A9D18AB15966F626486373BB0641FA98E0564A979F6A5F6A9438A4F10E4D2735B2954289D027B0774EF850FD92357D683CC0479B3939FBEC5B5BD809DD441F996005F184A9375928F183D09A56BAC56D4281352DE6873BA319ECC02A4FA2FB1F93A7B757A2BFEA72EE2E2374DC15D81B8628ABD863B241175D934493A9475615F8ADAF2FD54B95EE5A99E0289F99375E7F6972A6B7F3CC42D68DA338AE440BCE56C30E14735884F8CE63CB30F517A501CCF2D7B516ADD806C122875A44645125C9D53F459B0350571F88548FFA8E655DE8E79CFF6AD5A49608A917C3AFA48123F2C5BE5B758DE968F2428ABB44E0AFD9E637FEC58744EB8830B5D2846B4299A9439870A9674C95E6AD2344555DD54CDB2E8306494DC5BB626F25A70A74978C3698E89090BBDE5CEC804C8A42A75BADD8C0471CF7793192D4292B88C33915333766EBB10BAD0C224A7A7F7BDF99E48EF8E9E020A8CEF22149F33D9DDE28D66CFC2C2327355396B8E1EFEAEA9A7B8511C609B09AA512605B8D2105A265ED1235641AF665ABAA98A8838533082A80424F95A38BF05D3B86F392CFD2CEFC1A3E14F7156ADDCA1AB551FA0ED62C05F22A60EF01BCA302094ACFF7C18060FC92B759B138FA55E0325151478DFAA80B7EB51230CE61B473EF4DF26A4A0F1B6CFCDFF4B7E1AABA045A2F50B62F934FFCB51A07DDEC5DDB876E3A5CF3FFB00F820781DADDF65E258692FF8DAAE822AE4B40F11B5A9223EDD7BCEB1506314D03E8DA39D9DEDF90EDD0749A00DA34987284418D400398E9BBE05FBA6DE42E9A2093DAC1435BA7F0D981F4B3444E034D9129CF44A051E0DEAA1D9480CEB811E284B8E80428C5C141C8E2DF20E142064F602E727EC6B25209970287059D6FD2B8A2D5F64A9D647B04A895F6F35B77E1322231EFA071B4B87A038668A4C96AD7BFD53A98C274298150CEE4327E2D568FFFA7516F742EA8F23A986B731FB44AE8DB142449EA76888391A51E4963EE50E677A51DEFB246EBE31F240F4BF8BB266F184721CF13CD351C9703B56012C81749E3642F46236330FDE338171F931F87470530117B38344AA6EB4052E243CF1B3744A26B80022C9F29C35A035D74205DE9E6F92F2DFF5BEC4FE43172C38CF357E7958B40F0096E40355E10D725832ED85E04DFD59BB6B1C3849274EE4361FE3A9A7F878C4C7F61C8BC94E5DFC2E07FC4D275D4C1C78DD76F21D8BF51D22AD51A3DD3B7A447014D33C5A6637225D39B44E44718197C3B0E5223CF8D9AB2276F1F070BB25D24630BEB8E51FDD5DFFB3FAF7271794149DC26EF31DC0753ECDC84C27B436D64820DB55D8962F5A22B3F2E2B237A7636EAEB637470346BDAC1944D84F428140E26622AE9A8632DAC5196249CB7C9E83A6178EB905294C7ACF65EC1B60E463950DBE5F50BB5D8AFD57CB50937E16138834B5CCB2D78F0F41C6DDFC15738A9615ACE06FEF04C33962CA5638146B0358BB8B5FA5F70A10756D9D5423E4B045439FDFBB96C6D1AEE7DAACC6C34CFCACA5EAC2BC6AC71A65D143A7418DECADE6399D9324B100EE1B67E626B06CDB541CAF2B40C1CAF9E2E6B480CC84D249850E8B19A227599BC7F6AC8DA64DBDDEF69DD8898B12FB28FFDBC4FCC089079AA91E23D49F53793CA63A3E3BFABAD5A7E38519C42F7B57B8D32A6D1B640FC6063297487BF591540051F804E2CBDE535CE7290C969F3A31E19A1965F353CB24BB1D0A1A4E17CCD0E01BA8FE516CF1D2491DC0E688BAE3104CE55038C6817FA9504971D4AE17611DDDB1B779AF771741D2EFF7630D2B7E2CF1A821BF359A82A795586568AEC4B23080CE01F6D7D4C86E9495D359291501C5B210995057F1EBDFB89F5E77D5ABD7A63920881EE1204D8B0879A1117A4B46F3C04B14866AFB5108DCF327156FC0E845A74D947008D200C6A7045BA90AC8D2DFB4BE38CDF18EE3DD9080E0F1F6E48F5422BBEA4D1AFBA2091916054EC8E199CDF51E09EF251AF1918ABF6BBADB29DCAC43149A9486C7FDBEAD5DD8F3106E8D0C3BBC1BC380D268CD40610518BA5F66F20915BD55FDD57A00E19AC18DD841F28FC8260A321BD5C2006A987A00D8DF596EEBB13512FE552245FE37A952D2D355CA71DDF813BE42A33E28ABAB101B68389AED94613E1C746DB039C884BF13FABC15A89579117A37035CFF41875C156C0E72F6CD4D8EE90E5FEAEF624AC1AFA28FB007B08C29EB2F582B235A4C7C5F4D22848A2461A3AAB3C634BF5430D26236A74BBDE69937E088A75860E842BF431F4F2034BD0846EE4D96A0E87CB28287C91366098F8B9E7D5731826B4FE13154BEA161E6C89B75ACA0CB4975068F221B02A84229976DE48125E8C022A4E7B9871BB7779ECD95201B3D0D67741CC45627643752F9685D0C26303F7BE8A6A2AA083F56496CB6864265A1BA76A38424B0A1D176D55EFFE8ED55142E15100AC1C5B3A0EB98CD6637AE398652E255B22044555F76BA7C565AF3D823AFA454BFC8B8840028C3D88A10189BE33BA9E3C10104C872D4E8C355D5DC74B412ED8EC381652046A356B6E8C73A383A004232CFB7FB012E67E624F90F3766DFBCAFC448529C357E79ABBC1223206909E1C29D4CBC2163D725D16FC6D3A9E26F78EA1930441A0C9D9EFEF11BC2270FD7BD08A2E196DFC9C5D008625F39D46D7AB78E493308161284A4242C75F733EF8830A99B4114A9EDB21D1146569EA0C1BB74F84FB1BF30715859C78B8481D6E7166F01000B8FD273073FF873796E6C4C3FB8BE5CEE5A4E8940B52B2397A11DAA809AB4C2EAE07A69C1E6A9F0488136737D5F3C923C6781DB21EBF085F9A459B13030F4BFE1D9AB7C5AFAC460256075314B24C7E1525DEB854A969C866CC5549656CF60BDB271A835409EF027ECCC61CE725D5B5E3AA070A0FEB7218A1EEC1B4B12A13C973EE79E96830291D2FEEA3C6C20BB72781077378356AFA541182B47E271EF1229388279E4D56BD57233D74093F839B566CE8D2A24DA7519B8DC64025884D5BA3F7E34A5D61241053AAC01F8705871B51A83CCB83C1E805DDE689C25EAA681843C579905BD54392376C938B528437244F24EA8EA090201C883E1FA1F45C7CE73613A4BF29D7403C36DD5BA4DE7143FC877D1EDA919E2BE784A2679B117A6F931071FD9581BFA16EFF7C2DCC77A5BFF0DA301C64EF8D5934A9267ECB4540B963A9D3499D621E2DA3E10E68EAD3D40D026EADDBCBDE1966590F5FB3AF62837C686700A185A82D9EB6FBFA7D55E768935DD5E04EC2A820644B58F1CB00D4299E5F644F536732E2E3BD6F84EB4264BF4BDA6088D801E2E0B7BA67D3688BEB0D3AE73DE2153243F3E5AEE231A25FDBCB1EC07DB60D0E11DB417982965B1791C5EE12E3C60E8380C9916D96EADD23593951C2EAF951D9201EAE4B6595FCD4617C98BF54FC992C8D09BACF902E2CBF27A60E7E6BBD932984430F7DF29C8C3A98219BC3A904CA68B8BC7F7E23D61C2F9BA1E8F2CF94F6FD4042C31E6451E80D88DEA5AC5DC8600F98DE1361BAD46C486273CEDBA915183DCEF98B0A146246CB1D3A538F1F7EA36A7C9107E8D2C4F7CC4DD881AB1D0647DB6DC42B0032DDA19FC6E526B2A0B920E31FECE1F1F08602FAF9BEE8B5020DB144ECF3493F62C2565E83F76FD4BFF18A368E84B8CE4A34CFB7048EC2883C249736BAE5A32BF0AF67D7BB2C25BF3E0688BC4725DA99436C298F1E39EECA99118BA9B7ADDB48ADD15B681DFB3B74C4EDF1F3595C9AC7CE4EE3962D51FC4B1785D3F6A1EAAD2FFAE219E2EDA8E8260257E01B8506506D082C9364DCD52AC7B4481106223DCBA50976FAA9CAA3F461B3C06C5718B193298CF5336C8FB6A5F48CE385E10A9CE66EAEF9CC1930DD633C99221B82CAB6AB39291BA209AB7A9ED58F2A872DDF8D83CE42360DC4EABD452FFFDFE62E8C351F1311656F8D6A29A4BCBEB7D6760C621C7F50A7B8E9C9BD9F99A90D3250365D8D66A19390FB0DD476FA1FD7818956EF3C32301D8B199BC0A6A1617C62E124C49340412D6549944C9CDCC053A96F5E00150BEE5714CA9DCE9306DC2448A9B0364EC947E0896CFB2B8945E729E72FC683C6A9261217738EDB21CB9960751E918405A78370F325A93B1E06CBA3A5BF992D675243DA2EB5DED23A3A0633A7193254E88DE8805D2DD50A8354C8F646C81627FE417AA7737A12EE28E19EC92F2D8FE7FC116BBBE6976FE1F9B75440A407B3D903356037012F655449CF18CC0FCFC1D7946CFDFAA2195D5F787BD6D9CE5BBD40ADAE98F1042453FA0B0ED543F6E75DCF90229B614761879C27655B542971621F120FB36C9E52FA30CE455B29B584C4D3D0004A317AD04F611B3743FF54213F66388BC8BBBA2DD0DB54163197C3A3D36B64AF7669D79AABDBCA6E9A6F2D4E46FFDC1ECD89EF2982476922CB26AB1AD0B6A6714E9B211C850514B8E43D7539FE1F3CDDB1935979DCB34A98865D9FC093AEAC10A92C6E83DC8EB22602CCDCCDDFF0806BE63FC87DC64F9DBD1EFEAB372C1784C00B552A7E8B221C7A1020C87A7069963195CBD7186FB865D3AAFAA6F909C346CA464D3676221537BD5838352C2248B7C5F7B4FB73E1CB0D42CB4C94C3E075B3464CEBC2282E8EE6903FB9E47DFA311F3EBD866FBC0993B50875650508A676763CB62F5D4286754B6770040697D483A7D0543A3956B16976AA2D489E7AF556954550B801A1027479F7DD20257F3DE35113DFFA5F3BBCC7F4B7D160B6FF6D29879684447A259787CBB376F61EA620480AE3480BA37DED1A89CBDE9829CE27EFEDFCC746C847C69A1F83784C554593D34FFA2EDEEE5B254FDC4C8B41C0B70A44FFCC3BB17A704338C23767C9CDC966150D9E4F331227BB29AD41B60B8089D1874D4515BC5AA0719F2E4005AA84D39193580BCA913E578915899652EB107179C8E1EB9D5E5DBF21D82F8E8B9B3D44BFFF2DC77DF951B373EAA4737C7C78A12EB9DC43EE44D3BF5BD5051B44B1412D880512CA8D3E2B550BD030701DB89526F4743FCDC9C649D2CABB06A84E5C83A35AC12B11A26C166E86A60938179E7A617E5378C8559CEFB416B437A3ACB2FB1409470E9719137A6C3C9469B97A6087025EB35A4A718CEB695945241CD95202F05F84999EA0D814D99EE954400549FA3BD110F6AFA25B98A2E6AE702EEC185591D56E02749B58135462FDA5092FD117CA7311342EE4D85E62F835F6B32D77D643F384121D136E4C053FDA8801BD91D7DD629EA5C35C4916E88C16E2E85E522FEBFE639B07AF7A6819D59078FAC0EA78DB1E55065D62D4A78E8BC1977B872296B7D449EB356DF63268FB089803D7A1A924916A0AF50A0434EA9908FDE1E363226D944F9C6A0E0A46294A106197BF409789A37BDFA98F2B0771B4FA40B31F7C795C9F57446E2B4D9F70149A201275E9E5D9BC1C5E5DC0C1C5D8BEC7B7AE7B5BC36A23D780A41A53A501D89F6B5503C6386CA9BB0EE2E79C3420FC5EC2D14E781080EF23D8AE558E94CAFF45FAF4E2C137809806268BDBB38EFB86D532AE1EA547D3934E163A46D172CF46EA957598BAF62E0CE076964BA4CE065E1F80C85EDAB595BB92AED8F043600F9D722FAAB9ED1A069E9089D33A03654226077EA7E1104275944F62B3C094BF96B3B199B1E6F40DDDC761D8A05049E41E466F6CB0DA14C03624169FC6CAE1687631DA1D1F21ABB192B759BBA246668C33162D95290AF170D0D0BB5D9887C43682041E07DD7DFB4CDB9877A14BE491F281AE268B01646C9538B79B1A6E874A0958A4A03338E83A5AA12EFA95A02A286BEB29E4E2911DDB233757EF17D89C7BD52E17CC73507D1B6691B8A8DC88A4ED28CF73B7E95C78212417F1B0544ECC124A0B823A8D52F7DFA313415AB242F214E8AC3DE3EBE7865768A41E6A2F202FA7EB6BEACF9D8D9965B35E9E70B4E0C5438221D083F6B87D35DA1FC726B8AA3D4183F53B78857535B92F349C691C61772FCBD7156D62B29D27E37044D346C99A4FC7BBD12B0F911A978E333693DF61A61EF20EEF52F905FD54204A09A00DC4EC66C77BCAC280693DBB290F735F07BE71ED115197332F62CA927E51944D4C44A701923D51504FB77089411FB4C4987BA5B59856E4B4C67FA319CB1A7AF0F37FDADED30BDBAC740944F5065DB3D27B96ACF84188CC26227B0C6EEAC65A93AC76E7F5F1305A4474E73E647D062FD3ED8DDF26AD2667DB74CC0E2E4F4F94B26EC1FC3530A05F5BBC591FA96341F331A95CBD7E78C954A8AC1896518C179E9390A2A67037D82FAB0C58EF02CF14F30A1D9B45EEE325541432330E604C6CB4AC5CEFBD574C10CCEE4AA1A4CDDE87DCBB78E2BD40C3FA824EFAF28103C77A4CB026CD89ACCF6CEDDBDC09E866734F07B337D6DA991CDA7AE59B8DC439EBA8F73307181CE53A1491537BDA1B3EE01EDBBE2C6DACBFAD54C942B3C4C161BF68B5F747C9844F0D3320E39587EDE51D2EAA5DEE83A2A19F3FFC8C67'
			context:   '68F5D7FEC146227D50B240882B55E073604E69320888C089D08886E44B3861DE9C2316393BE07861BC6402600A1C6D1D4AE182E3FFB0297F2F13DF3AA8DEE152124AA499732A55E33168E23208EF9CAFC22EC32D8B742940BC8A6390C3A9CA9F960A4FA7CC304C0D0F0D5829F0E60992A4A2E3727E785D62F270C9C03864F08991D31811824152A6A142A6E8D71CB1864A9CF4B4335C73AF1CD2E81ED7ED50B5F62F45A26C532F985717CEF1277934DB8FA0AD8819E7B9D7768565B1D9AABE7033'
			hashalg:   'none'
			signature: 'D76AC1E3D253E976EA65A2AD15C0D8BB467FFE9DF2DC2CE12E212BB9D9203381BCE73A1A4A7D8E4941B98576CEB8BAEC95CFBF7FCB156655532C6EB2BEBE453B22E6834FF640137DECDF4E5BEF6058DCC914801FFD921E3BB5774630F0FD4611834D9C02487EA69D9280C4A3F288E02C0B95D4461220575EDCB8CEEB342F28873E2FE1EEF7EA8CAFB8E430D5799803ECBEB00E8693550237961C03BBE71F0EC256A5CD9EA48C75F077E2619309FD35BCD4351A5BC90B04D4B5930D1EA2C7686407FAFA6070D42B15A38919F66CA4C47EB803D3F4046BBF5E8C078A8A3FA497C39B3215EA91480B945FBD2CFD129F327E960E065941AC55FF656B78D25A61E003AD10A5DE41E83EB7D2507ED364D8B93B0E49DE025D4E0691CAD2A031445B6EDDB2FF45C3DA1853D775C64A7E5FA861F64C4F8D018002C80F83E2D859F37EB3144F275FE8F714548B67DC1884B22EA3FE44772F49746DBC0E1B73B5A8C82BC702B65A2832D7FDF81B1CD019B7A3E86E7A7678F10977E0FFBD0373A45E2FF7221CCED20F1433DADB4821B07547621BA69C9767D3436F4261BA215CC0EB23F18BE88FAD3278FD999BC39AE0A9CA39EEE27C083BA9C2D4E7289EDA9E8D874E14C31C45D50C3E9AB870FA8CD651621D9570D497B3488212C47942B5F152CACDF0A0246D66D97C8EA35749722D0BFA5C9D56097DDB9DE2B417E016EDB65C805B246AFEA2AB8011FBAE848D94916257FFE5F9937A2305918F0077516B4B780565FC5C5AEC14ABE04AF0F35468F4952F67A3678B57255EDFD4652FC8AB16201AF336EB238CC2414017EDA66614AB75ECFC38E5D2B8690F77F3B4A8DE98F7722053B6FC2BC842030913719850129C99A1D8F2CAD1560026B79B1DC7E7B186E64F59A434DD16691FB6A081DC5700C79FABE60B8BA20B11B8283CF48CC0583AC8C675119243978C42F81CCB97A1035948977D3C0DAA74B5F130C50FE09F1788A781F20FB40632D507B492B4F7B3C27DC9780309344FD6131610EA4FBC3ADC73B2E02B6FE214B7D9665BA91D8CC037B06B57A6BD3CA8496692864D448663D197ED80C3DDF301CBB41F1C6FC93B01B4EB47D67C3FA934256FB4C31A851C97A03E61216946943FDE10E1DAFAD7BBB878927D5E489A6F5A32E434AF84DF3F9AB25F63FD203A1CAB3A828B3D6AF3FBC25E620379401025F86BD7B40A6B8F44C304744A9AB2E3347F5F8DFB5FFE821A865EF66FA8001E4D8EA36EC63460E6B028FB8C49E86B9217F5CC11BB48F23AB124BCFB7F3E9AA209515DE569D43495054644AC3222BD87283BCABCD9DC20425B83A8549DBA19B34C74DE6EF9C6BEAA1B00F9F0EE50EAAF18EC2D9874C6BC46EC457BB12071E24503E78494F555982A2F12A88FB34315474791FFC2F1E173ECDEFFF5FA81E3B817624BA54F32E3C53B7D55DC1991F0398718C86BD465026DF7ACEC2839FCA48750FB68904409EA509312E7D2F17EC0B53F3CA572BFB4163DD1D83986EF107A3619E4B79355893AB93C4FC3BEAF5A0B87DC4E35E2895CBFB037C5AE85C4D1A3DB9F546C659499DB5D5EC91903CBA82E755388009C290AA35DF1A9BE6BDF2FE7D81D46B68940C9C0E6BC8376724ECFEC99420C20202414730ED7BF7A205DFE06220A27D107C94C7AC734ECB34AF727714FB31494B7E1E1552463B58802B47EB389C0FBCBF6B699492610767CAF2F5D92AA6C627AE92216960AC145D198752C499B14935D5DF1D3890F2304ADE9FA6F83BDCDD0593FA8270792EDCC838B038AADB7E3ADDC8DFAE8672D08DBC785FDD311B10709A1196D4DF0024843064E8DAC32C6034BDE7BCCD0147D64625887D37A6FE70C84DDE660820466F9646424AD253D2CC686ACBB172383EA6A9672D3260AE0F3F5AB0306168393839F0A273DC206C4E366DA0CD4E598E26F054B5F296F4C9907D66504A5EC25F6EE065994A39610507806FB45BB117D6BC12181676395A8E9F6FA7ED938F7CBFEA6B249FE18797AC45AC56DF5A1170123F210540AC15F98EDA298F91FA33962CC4A4B10956E26AC7474FEF4F721BA39BCA8D7E42D773DFC4981B9A3A8EAB5308F64DBB0DA7C5E1D137AE9B3DAE1FA3FE4F2496F4DB478B9CC0739741B43C49AB174E2DE40ED59027D3C7154305B4446A97D48CD0CA8D49F9F2FC04F212D8F370B0286CB817BD15AD7006303B51575825910675A152B7BA625F1EB56E5CA081BF5FA596C79EF027DDF99FA88100AA1EF61ADABD91F3E144B5BDA512E8D1ECB6D516FDC94192D36B7CCD923A6E64AF796C13C952F946F69C54DA3E6115C840CB2691ED9D23A84C724453635DAA346F3C089C691D5282FB16F825D854FDF51F08DF3F5C50094AE29B0BFDE44A394AA4F8AAE264EFA1E2DB54CE452377D4B4990C30A57C43446B08B3A90BA69544320F06E1A3340A22BDF88C6DFCD2A179C1BEF5535B8601D934C3141D4D8123AB4A7726AC433912028122F6020DDFF0F3E532D936B1598601311E039458E2E77352588ABFEFB03B09290220A84F85DA2C392C624B8DEAA596044D3C4D13E21DAF50488044184E7A490CA870F382802BCE8BED7623EFAFF07AF25BDECD9D5A9B0007D1107389A60EDD8583A8D66B2FBF11ECCF1114B946F71830EB1CFEB61A82B9D0A02A0C978BC5CB35D231C01947642804077D6CC72E34B48DAA8AF0FEA8F13A0D0E69C427B85B22DD64232C1BD28FBE3D3FFAFC60F95BCBFD6A021239660313E614F2B9A49CCDF2C427510E7BD1848E881ACDD8E3581A7538651D51B92B19CFD7175E81BD7E1145A5ADD20126979C6A3BBBA69C6EDC16235C1C56D2123A12B0287B45A9004596760066B0B97494225F6A311E6E16879B5A601456921F54439FBA0813CD4EE8EB8D3713EEF760685470A1E18A24D35E45264CA4B96B44A8A8E68CC4CF7588E74D28FB727F8A23CA187E0271903BCF88212615E6BFE867313F4575DEBD931397DB12EB5B7F7B02E3FC0337388326A154C1621A4727917B7C44A87A6DC7DB83C5ADE18050DD01B62DD1D58980CF8F3F14094FA2BA7A1A0CCC837D0C9F4C3E9228EAACCD8397AA313428BF91C2B97C0D39C82C65935904A460E92DB82DCB763C88DC2383B8DA923234C2A2819E81C8B4018C1AD8FE4636CDD8997F7AAB76F8D6656392D23728BF9512792A1D0BAFE039F7138D711D5CA8DC997C8B1D6159239FE963DF78CE1FE99493CAAC8D3040562B655C8B52130B03DDA780767BAF28FEB131369FC41FC01FA267BFBA2AB540E91EEA54DCD10A1B6D84114D4589C93727C3AB2576D73ABB98BD26FB287897EDC7A512EA0497FA9A82D958EA2BB3FA0B6E10C37C3261D14467063FE446A2EDC40753BAA871C4A19F9A7708C06C8B0790870F11A0B4E3C51D0C9B15183277AC906CB271A34D1A0134664A52780CFCF6FE4EB65FEED34BE5DFCEE46171D1E3AFF5E84B28120F8BD0DF74F36D49B0464F5A50DFE5EB736652CEEE16B37699DDBF92716CA48896198984E8DD019CF6073A5B7CCEC700DC5013A3EAEF8AC4AABFBAD9F41A1A24F867D405F513D829B5F52F0E24D280D334323CFEB107CD0ECA3B87CED44E135E441D765DF737026EF69DE43E5E795DBFBDFF69F197EC5DAAD40A0A702A4EA48E94FF33757367DD71B0093DC65F1CED71AB06C8E424852430A6A37C9B980537C3C6E08326D746A0660C067DA7BF8452B76109E7F8D329B6CA9317A7F8DB169C42E8BBAF753B2A9A5D091C9842D875BBD901FE1725DAC3C76CD1F23032C2E5D86D804867E001A9D2C07A20690EEA4AA68282E349E9675E8A39B2E3A74D5C08880238E1E5DD3EEFAAB8EA9BF6F6DFA1790D12B5287F27E57A7C5A0B59762D58170D24A9890C1429CAD8F2DDE45FF50895C432AA60ECE808985AE99F38AFC0D82C9D7AB687964818D86E1025A368AB72E262F73EB84505FCDEA1C8B2458CB588EEF0E7F93F8D4F903ECFD79AB6610A7E090235BAC3D937335FE30856F796D5165820A9F6BDD5A0E4070D82293E50D4BBB0394C63BE9DD5C1492F028851C0045E96939F07E1CED8DDE08A7F6AF47CBC937A28D59D97B1BF88C4732339D6398E2D81C751F33BFBCBC768DCDE34418D8955E31FD01527C4DE7F486005377E3E2672E93B1D3882AA9F5FFBF57E4CB0E38008011078224A38E6C6E9D00C1873CE12FC1ED912061D1D04D42BC3463A17B01DA12E3E05DDCACF78A5050DB4C31E849A2ED3CFCC5226796E4141F76AAAF81AC5349A610B4BCC2BEF0BB7160542ACBE91B6090FFA4E225C9558C3920E5BE0C68F5E8F276B6910A2212BC4C7CEFB4048BC6A57A50C24F858AEAC9A8E041FA06F5928034CF958F0470F8DDE87B521CC065825395C83EC876C3AD0F365200A8C5D20B29E6440099288684988BF8D0B9AEF4737BA073FA19C2F33253EB30AE343DE6316487B16E162531938F99DF3EEDCAAC845B88FCEFDC066FB20B92A309C16814A9BFA06A83976ECD58F684B279FDAC8617DC993920FC463A33FF3F9331E37FF4469AF22EB1108643698600E52007EC738CD737A3251913B72F6ECB7CA7259B50E952E135D09EF6F743A1479D8C2813EE38AD5F5A053375DBFA55117424194B4AD53410A12A4ABBB33AF6C846AF7B75F774260CE6F29A92583B958449927206E004AF052ACDA829DA7096A0EC1B7947240A7DBCC1F6E64A5DE903CB8E029FFFAA64F07C963AFE0C504FEAB16A261FE02781C90B9EA5FADBCC189CD7B51E22F0D30568C986164D6210AD2B6022ACB036D6A6123DA4C5FE815A2E5133343159F3E574DC16FE8433AEBEC782305CE2649574B9CBDA9F559DA4FC6947E4CECD9324DE65947D4037A021A3BA01965E14DDC76779CA7AF10552C4040D3B759674F1F329BF8D6A7B1CFD7D088D0CDEF7C428C79D2D81440F87A51A44A8561EE80AB2684254C0F14A2286ED93B52ECCA16CECCF5E53C061DE597D062A74C47BD186774B685213156E0DB513C118BDE60C69A8D4C03A545C960388EBC7AF702C639E159956D955DA6458079821176677868A840A84AE89EA34E241DC919C3278F84FBB32D730E8918C5129412D2D05E89D3555C981E70FFE9E3DA9B4CEB15E06FC05F6FA3287CB7D30C7A4032EF36177CE93187490A0C06184A5A218BBF97E62C2EEF3F11F6DC7818617C25AD187CACB7D4E170C265E4EE29BD504391052CF730633AD099D7CCB03D8093E92A02B9CD6299346602A79C2DAE2F596A4926B65DA92051B3688B02F7697AAC2A8F924FF5A8FAF8DC5E1DB9842B8F76C3FFA05C9CA81AB516C1C774CC6088EDDDCD846D21A4226D9265C8C4C9298C403807CE540C237F9B38F0720AF29E1678132D50A7CB882F1CBB73144AF2F01AD8FCB7018DC94CC7EF6E1747B75F68476800F32457CD555F07A7C91B9746D6D8BD065BF4D1230B7E83F88F2B9FBDAB4862FB5358B36E85B94B7541E051E4CF85EA2C27AC22C2975531F20F740511E6C6CB2314C5B29C970D86ED9F6E268B0C5817A81102CA2292EA2EC18F3E68152E4ECE856022AC42A770C32A923902E1D278B93C28825582A0856FAD683593EF76783E1EC3432E8C02CEC0BE24E0BBB9A70C9A00CDC0A5DBAAB43082743EF18B57B693E21321294DE73DFED23F054A5026C81A9FD6B87579E6873A0F91B4EFF20790B39367DA5492DD33C2850EBC658882E2F5BBA0722B4B1D076ADC629820FE3C8297CC7592244B6911ADEACA8204A582A840F5F7948B49846E92AB58DF0B5D039E4F040B6D90198BB0BA8BCE4B9D7B4EC88065FC89B1004B603AB9FBEFB3A524C1FA79997BBF7B8FF4DD5E0D898DB6225DA9ACD26DB93964C7BF2A76A737E47B82F22A9DEE6ACCAA36FAF6934CAEA4E79715D467AEDA51BC5AFF26A921A433E58726C0402468C52911733646E4BE6EFC904FBECC3D6C09F1D04AE563DCC8B44E36322205E15E5751754EF334143A6CB69E7F2E01095DB695E870ACB8BA21F73277F384B29095BA8A01187A6EA1DA9CCE4D07B28F869A78E0A667E5ABF788A7C02F954AA78F1BB2A6B4CD4D0CEA89A37DE366140670275B2F5DAEECD03E6059EBE5EBA94E10C78053CCE82CFEA7BE6592020EB96943000BA29BE0D9205F79985A05F4D8FD9F3478E8AE4980D3CDBB89F261D87DBF9F746C9CD9087B1AE24535165802F7DCE5CDEB49F6DF9D5BC87972D46355ACAAA540FFD1A2B85DB582F439E84461187523D6081C0552A387BBCF965DD96BEB22CD87C15E93D8B184787B0EF20030EB874AD0E94669ABBAB6A31ABBE0243EA4D5606A1E4675C38346C247A0276DF7B76E82944ACA90465A141FC4E1431D7EB7AE726ED65D90775D5B9A222D48038C76A86CA8237B2E620BE1279655617FC4E7AB9F3E719719CA632BEA24FF903B9DAC40C7CE991ED7F6D2302713B09500B2365CE2A7AFCE02B14FC8855D6BC9016CA28DB9382857B62C67697E122356860D776873A6E7D9E718ADA21DCC7F829863AA2647D5655E6676912FE9AD0B021E66C25D01BE3F4E0A3F2867DBB74FE10E80A47FAC379CAEF09B31FAA0F73507ABE820E3FC8B6F06BF22C863B315FBAD3E3D25867957E14097EBA7929CBE14EB01EFE406675189A8B0F10D908BAF7AE33806F2AD9DFF46145AB8D21264261E749DC96B69CFF550840155CE9CCCCB6179553D47CDD431645B556531A08E2AF2D44B0E63FB0C12AC6B6FA4D917D4C5788DFEDA53AADBC6EF6F74A8B2B32E628ABE3397AEB2870E6DF22DB0BCCE0660BC98DB9D519D273900E6F4D4D155E966D5DA16AE0E6A7BDBC0629954A89515A50A81D63F5E45788282DDDD3367F9BD0312ED361B60CA0EB7CA04C8433554C7C81014967102E4FA0082646A5A0F5BE4F1AF0D5A4C1D921070D424BB84E293EC4F0B1E816A174F7305AD764CB3A97D914E845CFC0FB6D31D9747047BABC3E4A31E77C8D2127DF7A504DF2EB02B5EE26438F9E2E728967B778F6BB8B549BFD1E31C9F4D510755F075E1EA6A38C43F057DFC7756FF43D7CE6CA09FD3B8D443AE4375CB0486C14ACFD704636F09D476F6A001C04A6C522A8DFE9F21D845B7061CDDB713ADA100D8886C7262697E4C43AA5D489BBA3DCBE832027C6D42635EF55F9991717AE70CEAD1D93B8BF86889BF2EC555A1FA99070ADA87C9CB7EEFCC92E048DEEC3A4331897D12B194415CEBBA92E487586B8197BA88796AB66AE555206EF6DBB12F358CAC15431F081CD351F5BFA34BEA518E7C66BDAB398E663C61009BB0855F8534B1EA3220BBE0D4CDC79D76632E28E154B4B5D14F2FCDE5A999B996FA9A836F3527D776467D3E4983A1222BCB37789E2335879BF9F54786CC327009A3AB3DBF08660F7D991E8F6C7DA56D93F498447BC883D1F66F1714F728F3DA8693C1959F8737501A41B07B837F450D718B066C42EAED3F30BCF4948D16614B4D6FCE486083104B2C711231C62DF7F1C42A41F078AD64AEEB2CF4C7F4AAF5CA614E25DACDFB2B4D2D2433B2D3186012996DB965900EDF59AA5EAD817863A0B3B0E3FEDEC09291883A1127562C116CA17F2F7230F4D71C8FDA2A9C247260018997B240A46E34C1970AD7732FD0A9E5F6AAACAF5558A1F9B0D629BB1EE86FDAA2F80E148A6A783ECBE797F7C887347068ADA71C03343A4C7F77E9E1117BC200E44BBAF2AB20FA81C362072DD85BEE05E7B262A8040656982A873FA6C58FD091AE4A3633361A401DD2FF2C2FC7D06CF76D1E63EF0FAD4F38B2BADE822D46D7B4FD1D403B30C5ADB2D2C02299CDDB0D4502AF59D7B76F29FDD5E04287BB430B455631C724AFBDE9DCCDAF4F7E3E911462A0956E452FC118E612C48C068E1B78C961CE2E1E4FEE708D40649A5FB3D11CE3EAC83C5F48C7FFAF3977069ADFD8FE496592EE9CD42A7EE3A2D4F2BD5DB4EF15F63A6859BB69A8C628D3C4E1012DA4F2AAD45C46C9B6EF28D06A4D5E4F5DB793AA447F68C69A16E0123ED76969115F083DC93260F2CF5F178D0297929B57D35FE9C08F75F4A56AB2AE2E707D6BD95DE828C94028D261C1D9113F26A99BB4F0ECC0266512E5D19056D5AACB32F31CFFF4771FD6563A3C89D659D1D7C47C1CE22F3E0C7E419988CF907502AEF7D5D1BDA347B89588982B94247486C320D303582BE5C4FE19CDF7529212F26CEC65CAF677EC2C87A9DCF357F43213E4BE5DCB0DA84307E1DD70DFCA29AC2C5D975F02675B6C492835710567D71D79B30FB67145B9C5AC58DEC326B667AF3BE86D97E4724712182627530ABE19AE7C754BD9BD07529BB85487671174AF577366FFDEF2FB88618A42447227CD94E01EDFB94595472FD97AB548FB7C69FD849474B2FA5DBD405A562E3BA5E660C44F5ABB5530ACBA7D1B3548A6E35BAA49DC4EE98E8F280CF015642CB3138945A3B6EFA2C51653DDF7C4B4F4C96EB06454A0A217C01ECBE1B3BD0D1B97E7C4828F21F192C10909ECFBDB8E6A791D24AEA7DC846F22F52E6B646783DD94F4871B3F231812119A8AEC6EFE93F6488FFE15AB3E18D7EAF24FAEFB8A273774D23AD9E58D861D70F634BA112372FC0693AF70FCEB6091AE8C789AA9FF89A8F41F327B451B2805A875312CC0EB961BBB0FFCE7EA145CB77E46314787A71057278B49B4F2F9024D07FC6B3F852D4A7684EFF2CD216D24A78236EA61BF833D3D44C58AEC144C7FD41A9C0ECC1DB64D45658961BD469B44814AA3DC638D48CA8BBA29CAEFDF985EE4916FDF3E672AE165CB25BCCBA2B1999886FF424C5F39079B0F619249433574B27D964C75337DCD86D47AB240C10059F721914AA58682F95A12522215D277CEA2DB29F47C88F6EED7E869995887D896B1E0C018299D277B30C7F11F48E431BE84C77F8A1A378151D251F655F7018CF2816DFB47C66439BEBDD954C0F6F0E7D725B327DF7BACAE0C6496F07E8A5932CB7475E5BCD249CC20BBB48E9E4DB0BD10EEB4DA6872EF5F7835B1AA298B48A60BE6F4F9F992EB2CE8D620C3296E16261FFB81F88EC9241C8703E01CEB1F417079F77CB5A653ECC4036447A8865FD95DAD408FCDA5F9F1863366632DE05C498953786105654DF6BE6962CB7D609DDE36A924EE79ED40705D884082EA345854CCEB31078FA86BDDA6A85EA103FFB13C0887B874742AE173BB82F34EB61A7B6AB1D73A8C8067C97D02B117E0972ACBE6B9D35DF79347C82C3574AA49E11FA0706C9A0386DDE457EEF33F3D5AFAF167936CAC49011F230B4682638860B07965578B69D42CADF5C7AE249E0A9F9A9F3FAE3092C1AC650C804F8AFEFA2923957BA924CC5ED58ADE9BFF7060F5A999CB5D76D1889518163DCEDC058C217AE77C58B26FD0B528BA5A266A2847D54527AD212750E872D844CB9A3AC512996F3AB39E73CD9497CA859BDAA81EDABCF4A4C82BCD26E2E550CBF7D7C7CCC90FC9EA04FE2979E13738A7745EEBF87B279AAF3A95CBC4B76F0F929E2E8405512669CD8FDF7226054B0CE90E6D7DBE257FFC921BAC02F7341A4D806C197CD3544D2F10C19197E7E0C8E2288F3226A71F6F6026FFB5DED61E3E80C6688ED74642F54EA56C00C64C83D3137EC1B123A4AE133C6022122D41509242173506BCE0E39192278B6163280A700778B325170301F7E0C68C567D29A6599FBEEE7DFAF3B7DF5E9325B1997976E70D3FB5125EB38D871436C56C94D5B4D2BA38A9D0CA5C2303F66BDCD9D6DECFCBB19BFA1163D95FB8596464671858E32D36A7434E4FA177C0CB2EAF9A3A7BDF5FFCF530E0AE3E2A37EEF187535E6F99A10ADC342D567C1660F879A0F43037A604B1CA6531A8F4B054D94CD7104113579628631CFEA7E44337FDC9F82C482FC076ACAD9076AAEB801DA02B7255B81C02CA7318E4F97E5D5B57B4D20B887D476A88A6392379688B93A2A0BC31D2B1D4D36B9175173BF042A663032E1DDC0CC0A8DF8FBC59ECE5E5DB9AD58D0910386A250DC9ECD6FF19CE4540987E3851124E9396CA1957ED390D383E599E30D2F6C9FE5C5E719FF983659E896E25D6B5C4AEAA7A32855F34E7E9CA09BDF3B8EA8891E00AF58CB1E82D0B82DA0F4AAC0FEC2F8349AEF124471F7697E59490D303D1FBE0770F77C32320BF78F82145233CED054001AFF81A71A63B9900BC5198BCA321DD43127C5E86C8C4366AABDDC0987000E959EF368EBE603CD3FE24FE164695B3BB3DF9D261FB9A5891572E302ADB7A78EF05413FCD33ADA77EF4786C9544BCFB065183CA63422E6B2D07F85A68C1414E2FFDDD2302116F87CAAB4E9CD9A1191D19C6391D309E9B84BC40274B65C58264E04377E63B919A694D8492BC339531698AF1190FD7EBDD4D52B925381A7B2E4A9DBD8812F456E0B6A10D639849D2E5150A868CE310F0830D92F14A6990C5E3CFF3964F50D138078C60DEDD20A060496106EEAF5A45B6F5FECECF8C6B961284318BD7DB77F1202B066EDBAC34C53676133884EABCFC5FE57DE0E8BD7124F907F2F538C4ED9617D795CAB214E54EB3847E52929642FE6ED5F506EF88FB80CCC5034F8CF2FC3A76BEEF90FBC47A00D25B189E1D2F3A0DCCB27B4D1097D6ED0B7E4CFFB9F1C3698063EF31D9F4F7E58A5720199764E327726F22F6656B2F3E3BDD06184972E156E65E5A3C6201EBDA3E970485306A602C6909D550E9974AA6F1455F16AA57F526A4CEA926BD87671C2DB1B045B118CB66E3BFF45859DA539B212A20E382DC813C41B5B8A9DE4E5E89085F0B7745813C1560CE7885B0C89EA1B4AD9281C8780B1DF95A5B6AA1570EEBD73A05FCACBC3A99EF9210C05A9F84808973A0FC058DE75680041DED136934FB108D0F715A9E2EC2C713A5902D351752F6928A2DC448E51832D954EE58F1352094FFE9B62EF1DF17B104C4B021ADF43D6B67C898A5DD4B4DF1C05D0E1874C60D8D237AA75FF682463FB6CC64AAB5BE229D1DDC0F8C1EADB511AAF114F0B715856F207F6E9B81259CE67F7169730D51BB972C7F71183EF2B5CCA193631254DE64AFD62DC2913250DD2B1155740104CC954C1C29D4F36A43749E11C29383B605A03471EE57380B9359946F2CDB4D6CDBA52A6F90DEA3241F02640EC52BFE1C265B118150E868BA6F50312FFB9FB6979BF553AD3404FA6D6D36A4205BC69F97F9D07EC776E0A5E1F537497E947E192B46B66F1DBE50D65C3B7E8D85A1F140F85A472A59EAB2D3A23D3F6276DE2B765E49FECFA568218FF6043C170DF84C4B00E873E0FC08B2CD5DE2AA7B4DDE78B8BB2E9D709A941C3DA41D7D9166400EF0042DF7BB9A50F510963014F19EC4C73D3E99F4BF2997B2B41E201C93BA0F4218A536999DCFD51DB0E26326090AC7CA391D5097787A8D32BADD5E9B09CE2C94ED8685ABE763378B53B0D15628163DCA2BC9F3251018A96EE553044FC991981016BE2DCCC354204A79561735993316D5E2E0530D61940CD9F22DB42DEEE489B077857075DB2B9CFBAA9A4283B1DA8D8B045506233754762B85CB2145DC883DE984D0475283D74AA06A6B5A79305A2FB516EAB8F633F16D25CC0B0CE43A156CEF1F959BB57A440ACE627372F336F1D530D574CDA578FD792425D72F1AA7FFC0F5B4CC613A65EB8B96566A680D0284CB0796809B7059DC01F2C42A39EF1538BBEFB61978F560C7767BB95032493861B4AD56159702382B1E8A267587C1145E1F1E26C61AABB3B3FE43A757E24E9F3615D2E7E30ACBA557FC3EB4077710D4471F48258198BA85AABEBD80F68EA3C06B4F0C95AD47BED8B89AC625B84EDE795BF73C0D07FF99E8EB8A493AD5FA15FF5E06F6AA5DC02F797F37669EBDFF79B041E90F211DEC7089D72B9F457C1EF83FAAD0510D869C3F01845CD7C49B017D85A02D78FF8FC55F29813F59611A6638C6681E1F823668B9EC8E75CC42248DB0759042D52803531F25391A66988B8F4B387E3B006EACA2C9CA43C0D702F1658358CBEFEF112F1BC98A13D1F78EDA58BF057B44B5B4C44C325496E6AADF282A615F5FBED46646F42A1A15026C020F7FE80A606483AB58407FED26A86A62D52C56FD18419A9A1E90E2E30438470D5AF8EE86D1A54C6BCCEDD383DCEB909E8049E73336AE349FA06339CB364C2A5B204E01F592A1A5B36C565D9693CDD711A71EFC79E66569FF9886E8907765ECCC8E8EE2064D07BE52BFDBBF3B53E65EB843FA82A96C03FAC90C57567040BE9A96590314F2972106739CB35B7E4C3C334B7D92AB7437A12B195F757285A60AB0F435DEDE98CCD97C4553EE375DB90378BF65350286AEA30617557A9AC961AB7DC88BB906EFB44A70E6E47362A062490BA57B78D114AA829B3A99EEBFBD6E3E203CCAA03EFC09E09345A37DABD8CECF65E9D60E3D2BFE12FF1901412EA09A14864BBF8D738976BE4AC764E13CFA430BE7D1BA276313D36B1EDA022B0A63F2A584DF6903E5644075236501709D2DB78A52F6E64A27CC5F322F3B86FAEE2EC0E8459C914454F287A52B7256BAE97BDAA986120DE527718B71519D82E1B7854C09D080AEFFF50168AD95BA487A5C5061F36FE56AAF3BBC48475E7CBFB33F0155D227ECCC3F634D1A6255D9ABE9A1A3191E52BD5EC22301FC926BEBEE31D31A5A529EC327D16BA85BB0FCA071C60EFEB4513CE66FECF5016FFEB2F13217803CC8573BB51162372EF8657CB91D1A2DFD75EDB9FC18EA8502880DE66F1E8ED749055F91ED9866E893BBB3D7928501F90021035E4F0C9FEE374047AAB324E42E17FCEE9B8581F5DCF783EC5254E510BEFF73A5F8637F881E3405BE6E9F33B7F5E76D847A4A627B8253EB0ED39A4DD34304E03B01C5CD0323E90178C4577F61734ABBB8277C272A369316EAB9611D99699EE3CC171442DF4FDE7A0DA05214FEDB675545E0CACD595DF61AA40E7752B601BAF5D7A9B0AEAC2A3E7D103E612529D0CE47EDCDFF4C09E752A17DA44F14290E8E2F116CAFB78D4A7BA3CF467D99980D3B379DE747D78B74B563129DC7EB099F5E4BA6FB859707FBF9F1D3DE17648FEBB6B68986CAA46C4066276B447DDCB9D6E4EC5C881F300D2431410685C4AAC052A1194385D16C1D8108CB88DC280DF0CFFD0637EB577E9A4D3FDCC847BC1ADAAD6360D1E80947D91BEF5FF6BFAC25DDF578FA6ADEA4ED57FC9E9BDB1E130F71CBA29920F0D1CB03EF702F1A0AEB144C54A1460BEEFA0FAC331BEA285AED093EF1D6387DDFA292BDD43EAC87630DBB51BE16711DB67617AAE70A99AF957349035113C63F1CA721EFFEAB1B24271990436C1E94663D7D88D14DD2492973A02F90CBAA0A7A23541BD338A75F4B550B69783B4B4C061014DA6A5C307965027444FB53D029DC8D661DED0B8C279A07D986AB42DE37598D6A2E103E91DCF837BAB39018193AB6C1E694CCD3EB97CFDACF04EACDD04F9A2E343626D74910164C00B19FB1C38FE6D5EE7D25247DE4BB91246E2D3EB05EA74D9AEDF4AE405C59B30C6D2A24A3AAC3EEA7B989C0A557237545BE57022D754B784AD4E0BE81FFF4AEDF115B27B3C55BFF8FD269BC4F53750D92DFD48B3D4D51978E1135D22344160727693D6E62F065FF48E40A1149E452EA5FCF93DE43EC53A42640779BC43C16AE94E120060C9352D8879E4B2956CAA25F0AC13112AEAD12B025F90FF3C03DE09DFFC4F04A9FA3CE75E96AC7919D872FDF587E77A6F6BA301BF94FA0FA94F6F219C0284EBF429A893AEB7803B91DC3558BC30C7ADF2EEACA7410C9AB77F4CDF7DAD2773FDB9D51E4F01C254D5DF34B8B1533306230E5F0FFCAFD8AACC493F6241DA8F1EDA2A897CE069BC0049B2E0264D49A62D2E3B834D184A99F16956F8E7098D2C30213B71787D24BF96F0BDCC4677892C9A97A4E845C47472FB079B22CA5C5546FDD9F3042040EE3BFF07944E2D0C46B07FE4623F559727CC912ACFB0710E3923FB24E345CBFDB0E831C599870E5B1E10752961469148C7F6444F873F83BDE8A7F11E8530DD9F0EA28806BA27D400BCF33D05B92DF8328538401E270C6CA323F33287EC7B6F236631AC3AAA74C4664705ACFEE78C05003FD7C7053BF2B072E303EDB236A5DD2006B92236F069EA0AD31C4C8B877099906FE4EBE8C41C4255674146C4786A58358FC1DB56A297429E454447AF968C55E7993D4893794D44D1E4A65F0EADB85BA590B32AA7F654AE19EBD6A1D493318E25A981C83AFE628114FE320CC670A9594232D19C5CAED6D89A4D5D343FBFD88633B25504A03ECECEBC4D1C2BB2130E290AE03275D3F9C3322BBF8FBBA00CE1C10B96E3D88CBEBC30E3601F5C7DB22616D7828EA44BA164EB1DF3DD3D331B494CB23D5DE421FF4F36C727F03C4065F1164C74E5861397955BF1865A93B8FDB7056587D07F0BE2A17462234A4A6786D28C9E046311C17A56CA4B30966B1662D0D9679D85382656DFE197C70523503961EFF449668C794DBA366C697C2F9FB93F762C4035CF68B462B98FA875901192F1914024A8604CCC9F5BF7C2EA77ADC6A5A640060C4944953C19A26BCAF988CD16D44EB3378DA5D340F72E9D510BC02A59E2FF3F02AA2E7B4CA7669A197999279D3578E1DEF43B75F1CE181B3AA8DB53C8371909CD3B7A18ACBF579E33887AFE84933C97B0F7869F2E813714AB6CB60FDCB67B0E03987EF3CE5858DF3D7C51E3FC96C51A51C1964DDF015EFCA8C349A93BC8A47A9BD03326E5AA3F60F1EF70D9B07BD49F86E73B17206880B1EABBBE36671512BC2C625330FD666E4A4BBDCBFFF3D9D86AD0C28F0A0CC03FE136DD84FDD866A925D6BB03F71446814E0B7F45718116CC06EAEDFFC92DD44A0B5FB6F200C08EEAE25C8567216F4FBA95072950D69EBC4983D440427ED299378643F75CF6AC694CC51EA1E619AC2A72749E0581DBF2EDEB000A894AC5039BB560430AFCC0979C8FEF762E6FF40C22421B40BCFF57A683130B90AE490BE588043278857261E744638F187B41A778339C0811BA5A80D40A9AE31CCF03C8DB4A7C159E5B9A78AAD93EAB11EB8E2EB3C9F089B6763A2B3526AC6424AFA8509C3D30937D1099756C682F661B635A7F3E0AF794D2C756F19E6D3EFE74ECAE39EA458BA938AACC7721C8E148875543F24B19B8346FB8A5436A888BBE41B90A395A2F1859D167788C97A67B9DBBF64DCE5FE0AA8E3CCF24B947C27479F33F447596F7F83F08E4FDA3E8D5C40E3152C51FB98434F4CA48B72B44BB1508350F54E3D0C9A5C5611C29964D407EA72A6A414CB487C89CD31F161EE4486E5509F4839D13662182ECF1F46BBC57BCD1CE3D34391C9943E6A1AEF3141834FC06AD25828AF23B103E6AC7047269FC3A80E82D69D216827329DB5F08D24854CBF2F80934BAC9269C53BB7333CFE91654CBA5A4127A63E20DFFB1058D0EDCA3E20D74278A778EB312033B37383D62F58082634960FB3E50E2764CF1101CFD111AD2449B0B8CABFC886036FA81162941BC3A4B60B450F527243E9A017D4AF4A3F7C817CB987484D1E5AE994495D0FE67A04F7A93C76B7F0F40995C3FA4CBCBE3716A7EC9E8DF4C8B8AD25FDF93FD9E69B39CA659765C3509096E7BE8FD16C4BD20EB06D2A189A6733695E5A05C411B03DDF99A18BC07FFEA1D22F24EE5F8720D39A1786E6E139190808B44B6943713FF7C5BFF90FCB0D87001CF09BE720DE97653D48A11BF84494A1A6055C73B879C381A8915E89493B8C17106ACF1F32BF0957D02D5B9E8AC38DEABB4C3AB1C10B3D1402EDF59C0DA330C8EF0CE2800A9EB2B1566DF1E0EE2999D27FE78399483FC077A45006A09CA2FD17F82DE6C7CCDDDAAF461AC7F298B31599E828BFE278AEA5B2C2567536BAB0F843D81C0296099E630D9E220913FA8527B35ECC2417C8F3FA087AF42641C2880F6393CEC68E48BDFC738FEA2F2F9EA0E01226319D96A169CCB63A8EB9A6E13FCF003A30587810C4A8C57D187F1A71B211E77E148C320F4946C341AFE0D73DF1A2C840E0DC11361F9C29612480EBF0ACA471D65F1ADEC96F4F60C186176A63AC84C463EDAF13A3A0860CC2F2BF79FB73FC61538C6151BC1AF89FAF28910F74988FA1FFB3DCEF08CD0F0F7B75325A3E2496CB1260D9E0DBB67DCD1A1B6256CD7C4632C70C65D3D706C52533E2FF5FDB232C374690DA3D4B6A05B6A6EEB8F01E1B0A6CFA0AA1418B571077C1AF6F26762B22956C31F725B7CBABAFCC32240B5B29CB6C50CCB6A3E617337A528D201E32EF6723A9017916B078546F64742329CB4BF16624D2EBB10C4592EA07BEC2DEA6135470E3B6C33487433F695227252DB50A5845130C86FBAB17B56E78C4BCF9D56FC93BE65E55B27639972C711755C1F992D861F404BE8F8563B3AE53F18A94D5D36B57EECB2AD9280AA4C0C0056696622FA6E15C27D99EAACAFB6841437AA21DB162F64AF9629765CF7BD6288247D9C4C9DFC5E109A34C85533EDACF975A5E61223A04E5068C137E5836233C9709C8BB2BD199678B71C66695A0EB55D7469CA8A6503844797211B8DBCE9E2FBFA4FAE55D55691E7C611D0CC5C03BAD970D68B9B1C0667D9DC487ADFCA3BF347987B3C2B4105B22FEF15A409631B9B0E3180E0ED84F3D6361D0DC0758208C7084E8086EE9F05EAE20A0742FF5CFC1A04F0A2204030979835B9812A517D3214D2BDD0B1B63C0CA0A63FF11FB7FA0891172E597203EAF36BA315887578917D3CEC0A5436B53F71FB4DD1F9B0E5CF4FFF50A238021CE7F80C72D31A2B74BD0F00EBC3C06822439A8A9B066E819E362E6EB8754AB737B30AB218370513E2A7F92A6A4FB359F9F08590EC03E45DA5D52405601134BB17C157CAB9B1DE165F1695A24B1B236521021487485D91B696E0804B79C085F9DFAD3EEE9B8691418B22C379FE446256E4B61F6B554D08F5367F6A929B30EA4C5342C84A34A214F0534CADA0F63A8E342800B575F5F448A5ABC81BF0E7D3F021FF04E059CF98AC70601B479B51DDAC8A433C77521F56B4DF8A0F9423829D2761B7779ECC5E3384007EAF612CEF90893DB74F109FA973F5BDA092D1ECCF22117791D4F1106BA5B78C8DCEE68886F1C2593798CFC6E0B37DF2A94FCC9E93990A29BF8E66CC558C8FAA8CF1F2A7180A34EAC3B88714EA80BF7A6283B03DFE94A9022AB1B9BBE821DF49730626360DF9C473E7A32AB55762C58FA72EBDDD17A65C1D29FE526FE3FC7AA5BAD29CCCA84E36B843E78B46189885EBE099B34E3D6BBE3AB0E0EC06174E4DF30D8A556F373B9A288A90C4518B4B1E83B20F19410CF0996584A3BBDAD0F93386A2D3DC2CB1221977240D9D09B44C29718AACC68D84F35C99B7F1AD4AB42D0030A49D148FBC7CC34DCB1CA32CF7F4CC99CAF2D654B67C843897F90D1A53A245E89DAF9A98509767CBA35FEA729BBF922D4C78F05DD1D44A4C863E412473A45C08C15B793A7656BEA19188C5591E80F7312BDA1715242F00060231952FA5B687EDA13BAEE686FDB93DBD8E4860B3D1C9769F31E6125F7C8FDA7B6484E24981A5C6D2479EF1EACFFC312375444172C451E47C920B077C71AF89DC3A5797FDD442B1C028F6D8EB808A2C3FFF2FC489DC45792DD89DA2474A6D28CA1CD491E1F0D348ACCEDC7B25F3E9065433752A355A69B3DAA0889AF9458C4FD3BEE7995DD1B49FF9B88226D93BC47FB71C29FB4A8B44CDA346F28FB19FBBD038DD65C881A99F6E56C25A4D1719BC27A55FAE3D1D93B87957C96BE26A59A4A64C9CE617D7BC2649B1A9FEBFA6D6036D8BB7AE56D759BAE37342A584DC4591FA86C8323F87079BE98D12F9BBAE15CBA5AAA490D8CC9464600A172877E765BE0D59F961159F4CD244F4E9DDE345A3F287EBF52F07485B815F2E25E1702BE99E659ED9E36145964528FE277F95DF34FA95450F22A7C64B1F56EB88405B70B831EA88E3D88B38BDF17AEE6EC4181D1B33F6B1461DC1E33EEDF61FE411CE5C70AC10DD15231463D743472C602DD2CC38246A115279A48BDDD53EDED1D76654B75CBE10767D94BC4A563A48328C717CA6D73E1300E08E5161101FB4AED1E829BD50DA68B76D368FE4BD058B717B1BA514D8769137542834B0A8532210FBCBCE9820F40434888CDE0EB26824A8A20FE3C56A856766E230E841CD7527D5162DC5863E02E5E01E09C253220E84517223ADFB51F5E762C6DB6BFC47FD4C8E772864E750E2145D0B9B202DDA789A3608C0637907C87C46A684660F4E7AAC09AC2D272ED169A519913D2EBFCDD82F85FE36112E4C25194DD6B8B47097E951CA975B6FDCA61585F30F70798951C265E02D227A441B9576C2B558166CB4A5AE3937818B99A9A1463133A9D35ED14E4D6CE40EED67D88602D2A2DD5329BA91D17607CC3A329A3B6CA5A4428543195123C2E20E1015563362E288DAE9B129E72CD2141208C9AE84B41071235122ADE1C02D5CF3766A5619CDC31975D5081D3F6E6B8D970C397EB0176F6FBC0424D2308074FD2287E1CBCBDFDA409B4B797C46ACEAE1F2EF3F9B33A773873A0DD6385F23FB84A99D8673A4BFE23A7094D54D627A8B33CA4BBE685B8208E13DAA730CC3618271C4E77868943904A6EDFF7225ED38D5A0343223ACA80929C4A38276D3610ABA6C2FB0A740FF1645B20E839F929AA4A547FF7CFBE86DF0CD5A483E88EF20099508DAC8FB04717072BC525C0A8F4653CFEAE7DA0598D7713A829738D0E0297761B66F26E0E2C7FF920D7664E91443026A11B6144DA02E5F5BF16E7559EA2BADF645FAD724FD8A8150C6801439039B7F6BB542921CD872EAB75F486D1F0E404DEFBC7AAE3182B4C91411075525724BD93A72AC81060EF25AB88DD3B9EF0032F59FA481C18B04279C043812AB7815B58F599BBEA825172B8FF6989C021260C02B7DA722D34E21CB3B3303F85C29C4157B6CF963FEB8E40BB673106F0F62668DA6651150523847FCD958A50DCEF0C37826DDE78A9D9B5E0B2135A504BC84786D369BEFB92250EFE21CB1899CC5ACD1824E3CC8A65F8A390EC6376CEEF2F032D0A77044E13E6E74A913568DBD38C7058F17386CD95A799C933B8FB51DBA9C8A8D0DB546D365A4B6A479B80C775291E4FA67779C35C10882609DC4AA1EFADF784C3E687C46A89886432517EE8E9977A55B98057E1ADCD708AB893EE554AFB05CC1586800275F2022C9D3334788D37F0E4652C3F579ADA5BAA6A1C37E45A8D97CF44E53AE1898D5E2CFBF8A86AAA29D36C811E7EF75194B3261EFEC0865BCECB34CE045AE90483C34364D77AEB78B080B5DC4F56F3231CD6095B18F1DCAFC93C0D167FEC6619624E27A2E130B94840784E96A591A66148A6BACB37272078A8DB2EA7B890A9592595A77BBEF79E6C11EB916BEEF5A9BAA7FD05C2CCFD0204D0870D67836F30CAF7100653845FF76956ED97443FA33986E3CADEAA284E2CDA8D41C391B5F8377F4F9B47DED5FFECB88F097C929BF4C1FF94CA56C9C6B91C734A3AB3F18474839A96B7DE2F85DA411082B24B89B6F61442D0D06E6532D7990F7F32CF3F8CE50602C193C1B0F2B6C9FB7288F40E636CA9399422D86E805769D3A606D65C275120F8695DF5844CEED0D03313E073FCD244069526F601DF9162510C3E2E5F53D8D4FD83BEA0462D08BFC8817D1DE0F3663AADFCEC1B5925567CF1F30C82663A29B00C161E486EABE8128FB7C0F5BE8B6609E9AE2404D0EB3DFE4E1E141669FABE4CFDEB91A966902CE9B66A7915210B955CA1906F0B2F2621982B375C4E13203CD49405044C6D0596281B5F430BF80D526B7D57AB5AE50BFB47F29C35FA41C33F09177325122D29B0E06B893AF7CA8119B92FEDBFBB162A8CB5A1ACC7E778C73C10EA1B9864793DD69169016CBFF172C2E730973F1EB285A87E3453C34BEB57528222B5EF41B8CF3C65B0C65DE48C1B370FD9240BC02283B298F2A5FAE2B98E9877D47F840493426468364F9805AC451FF72FFE3B80916D9E29B130F0A3CA0C334C4D4B924C6EE8563A22B1C3160C3F134D9140608045C9561D138F4B2C5C1343F2161DB2CB7CC48AD04A870273E925E9DA1E76514DB5BE487922E1A8968ADE5861A196F202F84C1D1BA5588D00428D5925302F2BDFB96C5B2FCA2D2BDA22CA67AD32D5AD2506FD0EE92FEE00B1AF3BC885610A38D9D26A4302EA041DDB8BFDECB1F43851A25100C633DDE919F8417A79AF166AC2E6E8DDA3FE9672186538467A50EE8CE8D0D21BF2779DA6A1A6139D2FCE1F017F26049D4F4E4F3D18BD3D8DE5E35C84AA8AB5C9A26F0F212FD10B5092119FF11D382EBFEBB08F1490553340E2C73DA25B3E0D50794AF1F25B3A8290619CBBCA14AF6EA8037CB0228A438CBEBB5EDFDC70C25BE3DDA483B62A15DA810A3360DC0734EA06C268923E8959871D5B03E01D1D6170430EEB840BD4BFB9954A1631FF247AF299E3C41F0ED97DEABA8C1B734B60FD8B8D1E2CF2FCEC061F75BD8831198B54AE6F48E1A3908EB59041B92DE2813CE59A9608311C571CB420926CEC2BC3853742F82253D8A348272971ADF7392B64F7605C03F80B7ACFA80C938EA672F29233B923F965B475A73ACB40A49E0EA4F194EFDEC3A414543EFB04DC6B0E18F8DCD87A0C35BAAE76ADDE609D9D378358041794645550719AC6EA4A847B16391F4BCED31DCD456CFD780477408E2A509052E9FD5C1841A4D66E42E70944177C69DB37A1FF779AC50D28672715B4C8C3DABF256137E89991A3B8B631FB86690B78C7D07DAA007AF12B4C30707036015CE08F0B2ED03FCE900DCF9D1D07A5809D9B4CE062756F76261A3BC3CB55F38A0553869ED3F38BDD54D386AA0667BAC4A7E47043830E7A086471A607DFB89E70E9EF532079CD60A93299F963F358DA1CFB5FDA0608265DC9078AF4FD6D0424C0CC003A3ED96E45E2DC933517389187A358F15A97A16E3FF22488119B9484C18C883A54A48B47411774F164C37BF2CE390BDF4C6AD89D7AF6692A7177D305536A80C63BF1B8F1168EF9A737F1BD1DBB48FF7BD860035E064F00D0B726F1CF485F54F252CB925C913562869B2EA7747AD056A6ED53BD93CE76123695DA2D220779B30F7B8DD04FB0B31AD85A306CEE07098581D9EBDFC301BC14BDB0264D487FBE3529C82F6F66FE83906D31314B36638CC1887B45E6FF789A8D974694D1AF9C2ADC3BF39160D8AD86CF1C1D36C69D4975EED1B414490CAAF7EC00EA9B4D3277E3B8BFFB8760CFE91A4F2271E29E8CEB14496346AD7EC6B4ACB22FFB498AE4581D426AD73156BFE84C08AD429513D147560C0935DFBD49157B101F439DA3822A71D4CE0C655D2F297E54C7F0F961DC896ADAD89748E8FE9E46555D6A90733797D5574F2C3466E673595D906B1416E7BB773ECCFB3A5211333B728A36ADE1A43AFEF4F24A9CAAC128F8834BF39D910ACCEDBF71F3DEBC95CA1B363EB5B6020E5E4F7ABA8C8F601F6BA5526147626F3DC457020D89EBE6641E68CB8903DB7C0BAC54FF6F0BA1D5B602A1C3BDF2577E8C693646AE1E76040B806D69B826F2BA23C1D65BA1AB133792920DF4A8261ECE34F9DCC44C21F9C1A523DAE05D8E16028368AF92D9594A9F42FCBFEDAA944794C59C4F2721402B518A538F47F3DFF65D7FADCB36ED04B3D5D4F875BE2849D5621CC9F532DC42DA1262F80042240E77DB2B302C02E7C01A2DC3B7ED43CA435996DEAB90524E0BC860884565EDC1BB89EF0F780EC21AAC8752CA6139342AFAEE852A100FC0DB17BE621136B17341609EC8929F5A14D968F2E314E71E67C85024BBD47F29FB12FC1EFDFD3C8C6D498CB9019F5B66EFDA4E15383D5F7735878305CEEE530ED85F729F31AFE0B1325EFF099EEBC9ACAC06395E5390321E41C752B36CD8BD8A4F5A6A90D96400667FA2C9BDAE7FDF2674BF85BCFB04D239099CA1A9540CD9F3C41A6F46E0863AA3D148E888074BC668ECCE49157D62D7B04A96A35559632BC354187402B8F95150CA29A799FF9748B3524AC3F60604E8E92F83184D5A55E5518CCA0634B3511802739FDD21E0DEA75D486B8DD3B66DFA3E9E6BB598F45B4F2F5238962A820A1ADA357C9BAAB8D7F5A8A683827CAD2956FD518FD29A69E2CF52092A34041214FBE7045756686B081E98DD3DA799E2B2EEFCC5DFA6EEE8F6D02AAAF709A367C1F1563C391EB4AD76499F1AD43231F0FDC730CB80F6377E377899D9F210B456B68635528C47A399D4CA5574A8C924D2FD0988F49D421013A7C0150BF2DD031F95EBA5CA74892F86C854B10C794BD1BD6F59EFEF2E5AED90EAF47F78A5EE1E9E1A4E20452CC42640E7BF8EFBC155ED58269AEA7230A7B7A644DE24DBF200EE4F347972D633B0971AD612882F505DE1A4AEF1588C4622A07A89E9C888303810939BC7E5EC75A10BCC494EBF3FB3D3BB428686A61AB8F46BEFC98E71D21E8B9401F2C1152DD2506E48B93BB52EB9A9D1637A3D732F9C9C5D731AAE478762332237899F62F6F2A2778FCE28504449240B2518DAB926761B6ADE43565728FDB64C4CFFE6CA07EE38E91B435FE7C4B960F18BFFC9B90E0D949AFD7EFD0CDF28E6E2E4F1055AF8764313078AE140D5DD7179EB5A617C574DA3A53857B060134E728F9EF9B295FE9A643B7F5B5B621E2A22DAA2A57757283630C5A7FE1D1A6A709912995C2B2AB6CEE087706DAEF958435B6726EC4D8DE4B308433F39F0C06226B560E9FFCA0E7C4A2C89DB7D1D970FFBF9DE2A6DAF4DC849EB87509C63B2410AEC515594DC2211942E11CB193134DB94A42932A97B71D42AF5C23559D5EE6C011EBFAD135E2A13762DDD04DF9A3785C396C07B74FB994B0DA6D6514AEB533FF9660EE6A82B0B99F608B9F788AE4A7883AAFB0A484C4DC742C399B094AAB1CB60CADC6C2AC5EC800B0722874D2AEDA7ED20B8DA1AE76C782D8ED3AA855A881E667B740284EBB3E952A4734DCC26C0FE96E0D3C12A2E263E19485EDC0E67BEE249E7478DB8E27495081FAA14849FA56D54FA55B6201D38F6F3F81F8F50B9606C5BABBBA82209A5449BA3CE24B68328E4B54DE27E4BFE5EB3A6F521AF2B189DFA373ABA88700C9FF83E11CF9082B418CFC5BF1D0EAA71208CE7CB5A78A16C4C17BE8916E52E47B82A1359F923A21400E17954A2AA8BBEFB6857BCBF2CAA3825C2C3FFDF6821FEF52FD654A3AA537783A330619638E7C9B2221D20E01F922C03251AB72BA15646F7058B8EB8B1FD52A05231F58317BB70E181052C72E4D0F1774AB078CC13184C164E70F91348EBFD5EC13B0E198453CFEDAB0F8C8BF148AF6B1B24D539FB299BBFBF23D10B8399725C1FCA8FF103D0B4CFFCC19D7225E79BD06DACA3BCCCAB4DF2DB8FF39F8781915325B7EB10593D22DD5AF1A5DB2C5AAE4C41A9E8D204D65783B85B46B3E7215721932018D2548691452227EFD8C0615967116E2826BD635A7E4371048BACDC64A7C756B71C7EBAE516844A90ED4D89AA7CE2768C197BCAF131E1AB599B745960815BF7EEFC381D7D4E893FC9322D352309D1CA398A550D8F1CF2D7F68D38CEFAB4CBE7CBA4021A5CF529FD9748ACE41D1BB1DD8573BF20AC94360B16B691297FBD9FE1F79C8A67DE51B61D0B06C96D8DC00C28E16247552A83C7FBA39F329E411BA0C3E052C1D5E9DBBBB50A6C82BF692B9E5587602FA9D980130EF280CE3C59B9AD04AA65B4D2A2511C45D8C1492671F44CB0C4F0B4B572F7DB2283662B737B5451CDD51769823379788697ECB6004D073F60DDB1CD48AAF976D6F3DD868012CF3F73BC0E1B38E75969B5D96623B856A0C290ED0398701CBF7582901C4921230362E82D8F08920B099AA78F6D19DC383138B212E5333268D8EC0540D062D0ACA41300CE9DE4DCB006F87AA39311D9C2B59337CC494CDB74CF144F5873C77521AE312443E791543343A284A25E0489F9C645C12A5943A8EBFE1853A45AFBBFB23FF3CCF6B9E89894F51A92B7301F8B1DF67A27F08B658387C9F1391D1BA7F0698D7BFCC841970F8D447008B70F4CB290DD26AFCEEE51D68FF8D12738B0AEA3E461180F3E50B3723D9E0F3533BA0C4E49827374158557832B1FB3E0632E13F0FB40A6E64773B69560FACCDC7802A6A114BDDF746425A889DFB93D5BD91401C099882BB83F1E217CE3D3CFB1B16B1272B8C14956B05C9238A91E425802FE9C34F48D02AB8C238817203B78E378CD00295EFBD5B5D796B15FE7B56859846B1CA6A93B2F2AEAB529DE4EBED201A5E4643F0E896043DE5A4D468B7DE9C1C9C4851B3B9D3BFDECF40A674D15A90A1953E15505D62CED3632D9465C5A353E27F7792A96CF0F3D90E12AD01AD8C79C5675F9B845D32B73FA46AEF0D'
		},
		SiggenCaseItem{
			tcid:      2
			deferred:  false
			sk:        '96933BBFBAA46828BD4CF83A8CD2419D7863D69CF3EAFC91E47B33CED9985459C58383F7579C26AFA6FE3E607DA0D047BEAE389D9E2F9FF17A69F4E0D7F4D829'
			pk:        'C58383F7579C26AFA6FE3E607DA0D047BEAE389D9E2F9FF17A69F4E0D7F4D829'
			message:   '2C'
			context:   'F7EAA19141FC80ED319A842837E68FF126DB762DFE49CD5BCF11D0E66EA37EF6F72C382E9938532645E881DE9DEE35DD60DF56CF74726F2F183AC99422C6D6B37822176CC4F0D17CAAEBA06E79E69699A5F3AD4556F7180E98FC1E6AB4FD11E556FAC53387DBD00D24ACC68D8108'
			hashalg:   'none'
			signature: 'FC58D5CAA886B6084B562DC42A3AD0CD1B73EE6903D652F91A3245EE263E9E63457DA72EFE9C36B2D7BFB7953E21EEA2A684789E530960D7BCB67266AF98DC5C1632B415BECEC0C5CB90568C41B54DD2392119B9405A2E7B4A1D453DCE06BA9C890F73F3447E446A1CADCCFAD98DC4015A082FC02325FA09403B55C25FE2B24B0B9B0143718F182B923E012E5D880C2FBC5378A29CE284E2DC494CBB269130FE831345BE28D2E7F09670A7828806FFAF643EDB53D0CD4DCBE08F97B000DD8B86556DD7BD156AF78D525652E9727AAFCCC9CD7634F219909FF598C920E156FFDEF46E827D7BA2108A6A5D8D45EDD243C1952158E99D2D5452291A4E6CF0ABD8840F77878B64060148921575870E68136C40A6DF881EC0F5F2EFEF2CAA33C425B3F8CFD02EC7BA87F8079758E3B650AD520DFECFBE76E72BDC88F349C592D327CA3AA76784FDC3A16A4A6C7462E5CC8791D92FB9CC0A8027F8DDBDFCC6459277ABCCD89025FB9CF25AC00951864F1B17B56E07F5F3E911FE44CAEA6541553474ADD407C03BE00AB4E541160BFF3608F8265BFA13CF0955C566ADE2C32F9339D4C8818148DCB9A6F49EAD1F71D4B711126BD3CD89C4A489839064274E35EAF7E7B77760091AE0F54E8D33F335B211AE73C221C79A8F31F29539112ABC7995CF7ADAA356228BA8AB46F3E8561D9DDEB69D21C3ABE3991E4D2EB7FEDBEA25E96DDBE20CFE950469CAAE2997897B8401C5FDDBFCB454D912DE30B8715316BF52A2B58EA918306243E88B23AA2EB0445AF6ECF827E84C4AE4F383CF338B1C63EA6B32D02BEEEE064B6193BF7BA3D4660DA0A5BB3FFC600C89777626FF833D523885208329554BFD179F67180D44DA5CD29AEFAD5C9F77D5A9C7CA9DC1310583A7B95579A5663F6F836B271BD6D8805CC878CE59889F23349F06EFA53CC22D198624E2D3432563E96EAC5957CBF6434001FA97E31131278C1C8C50093AA4A491E12EE697E9DD1A311E94825FDABDD32E33F19045CB42D8A532FDD99661A4A8CC568EDFEF558C0F9A9E26446A424FD3819F939C55C1EBA0CD4EED0F8FDCB67FFFA55C2057F10FE356A92012E39009BE0BE95556F7C50057BE2D75FDA0B95978086AE34596831479D189E96F5E57FA22D2ABD715B61130F73D7AC58E0096F862928DF9CE1865D6CF62E538D58490CE2BF34C37F346B7C498C9BC8609F4D6B5CC22D1C7611056ED7894E65312E4B573111BE2EB9092E482CB8D6E7E922A522D82882AADC2875BDC1AD0CE25A52299E3A3F70482FF4573BCBB7802C2442C1FDE350F71243F70E735C9BC6D0BBD1B6FFB86729D95C9AB76398F26039C6795C6E145CAEABC231C265D65114D116B473A0586D6213049FA0AD4B03CC854982A5ABFE0ED31AF65FD2DA994B109E55164435AE156E4AC57298601A41E984BBA7F94B9C560A6E2CEEE346A3C330D0B18983875B1BA5DF9901FD0C611D770DD9476D922720872182A495979EE9D98AE0237CF75BDC242AE42088A88F900124311259F20E4E7DB93A858CB5E3B868FFA7E0CF9CEAF37FC51F6EBEF127274F34C113BD0E124732E93FA883AEF53FC401C8570370A0A61896C57EF7714F5C374354F8014D4D025DB09D418D1F93A78255CBE899EB906B8A46B864C5339CA8A7C8062C56BE7DF799844266AC13D24508F61C4802B7C6D8E788C62DF076906A6ACFFFFDEBC16CEA745806607055919F74BA0787953C3401DDF831BADC9A0CCAE5E6A58BD0EB7040C1A8F31CFFBB9E99A877E28AE13CB26819B2EEB0F0DDCCE9950D62391475F5F792B9AB09C3F28922489309EB8C65FB1B901EFFA9E0C654AFBC6598CE781CB33375F49C929EC7680BE9A253A840DB11124104D56DB184B9140A27FAD8E74C86A3E2861D9225BA5D67FAF04F61FF9567BF1AC06CA47ED66EDBD0268199DD866E560C5C2591D6B900B20482637D4BD098F14B9C41C2299857D3391C1AF15D7FEE8E9465F8BB3448219CE65D310478303C738DBF9CCB9BF3F2C5332DA57C3D18F6DECC68A49A09AD16646E844F4FEF4E1B58066ED469502B61F60791FB9AE3DACE411F32CAD1032708FB54A7664F6B063D19505BAE03A444F38F49AB80B6789D975649D4C44C5829D58A084553BC7D64D8EE1E1FCBB3CEC71B89A4413BC850CFE80E6B5C125228D7140B25C4C9678ACDE76F635CC083AFB6A34934D153B3EFB898391EBDAD6470C219AB54D29F2DA7FC79631CF6E90E1015F60AD597128472096BDD9870F45F18853542FBC3B4E50D05323BCE381B3623AAF6BCB203C9B439A9C0DB3B567A85FB5ECCC3133FA3BCC6A47E3AF332A3C3D22C60E5686B36C140E51BF6C235B464181D669F65242230BD3D9FD55F82DAA66869D990A4DD88823613658C66814FC9299373B9F7F323AF08E41143220B9767E4E270B0AA7CE93604338E11BFFAB0482B050DBF9DE77C94AF055109969FF961315501C5DB6E867DEFBA1857DC0601974B2C796A13657C311D1C82AB1FD4E22C0F0B812DC9D9C6F7F4F9FF7E86AE3E36BBFC0A3CBEB9CCA5FB7FE4BC6AC08F6CFAE09DAE8E4FAF9C275E4B6E3794F80D422894BB8EB697960B2D588B5EA5210E0B3EC0AF31976A77B15CA00D487D5A3968ED4B52159F237ABF80BFAA75FA6ED869DC9009906BD3361989CF5264643CB75597E036571C22C451D78FC4FEB84A12949B3AC9E9C6E24D7882B7BC9C426A624447A0B0A1A757036DE42EC300811BDEFE296683ACF129C0B2BEAD7F07BE90F190FEDF4FAC9C91105E0451C5D4087B9C5E345558E3047CAE3D4C063970EE5DACE8C9E2C6D9A0FE6C47B948F6E154D6E893BEC0C88B2B0ACF96275B717FBB85FC6F5B39665050BDB8CA8456090083F8A4085BCA5956A4B4BC6A2D5B182E35F21F10BBC9CA840168571FD6D52B1BF1081A6C2CB4D51DD9AB51CAA763201C97166B2E962B154B78FF2822075151DD1FFAFB6DFCA23C93977AB248E78E353D9AE8DC197698B326E8D542F9F0AE02561C6FDFAA0FABB7F47422A0727100E3233ABCD009EFE7A53C55781161CC8D3B676E4B5DFD11582F0389B63696063F7B1562644EB2350726B4E17666F50A7863C53EC1E7445A1B28C688A0C4C08B7D9EF9864F348D737FF1ABB5D642FF5FD13218F95CF4D45050EBFD94D00E4CA94E06517A540DB5584200F7779AA2233D8F7DAD298E1336EEE51BE250EEF1300458D289B47D4D712DA3FAD1358582991378B334A25C09F7928F8BCF196A25B7270CBF04022C5FEE1EA10F0AC7FA6CC9159AA53AECD220652E53D435C9C6B164B1ECAE22416C68638FD9216775F89CACC8398888AC17B185C45BC6AE4A75F34561623CBEA79F7A23D7A39B4EF55EB57C79FABC6717B35A69D0B4A1F26861B8E8EC8DA9B6F0A9F7B20326E0E7E1A1D493790557D4AAA7A65B03C6870A030ED43E4155E8F08030F4CD16CD06F2EDE42DE49340D8F8954BAC29DC488973A77F80B868CEDECE89D0B082C885D6AC84CB4DA443DA874CD16373B65BCA862F7EE0161725CBF9743ECA7758DA8B5FCF653A7830D834591A95CED538D49E2EBEB2239E80EA04D9446B185EDD1A43013BD8A0A6518B60771CBECED6D3991811E8F527641EFDD05B4920A8D7A8A69159DFADAA6B923FDE8504245AAB7BA2DD785D3006AE99190B979C0D6D6C1FC0A369DC63FBB90648D35073813DD7FE0574D84472EAB43C002E8F9FE8E25F80A15435D9EAD5966DBD5B3BB2D9047ADD2EAD3FB437E2920B544B786E3CF291D0C9310015BB971481575C45989299134C5EE23BEB7AC7FF5364E16B1E0F53F32716C3C4AF2BE6B8F68B4172C500B99695F1D9A80CCB340B6AEB048FE21C721A2BED1E23A3A973CFDBE0FCDE341BDE4C3B5AF2B0B461539DFA62D4C56B51647289CB79F14932A16B8F2D1EF6F6FD210D63909D6D529CE4A4025E2EB5DD02FB8E06839024C72681F272B14F359D3F55B62BC2D05E23E9AEE64791F47739007A52A24DDDA30FA1D7494A711843D8A11FB41A10025D921B28986E474202ABFA5F480022EB15A488BF2F4A498EE0DA5AC99BA676669B854E7D7EF6973201A3E7F77AC16BE3699E0BA69F3871F10ABC36B367E867A8A20575998DAF4B2F265049AAE5D36DF3E2D3CB45803A649E87E28FEFE259AC8E506272D612146A652379DD24D45778B0797E12586AFE0E9F42CB454C7C532BD3FC5B4680C9B87417202705C21D0108075715CA04E2B8FE838FC43135D5DD99ACD65A2A1D48364E0044848A52F5880AC23F6FB5AE3439CE77EF659F93F067D2FE0C4432F3881DDEE7104BA6B9DB0EC14E5F0F6ABF6B9884DAF45CE70427E5B6BD5DA6D7A5C36665C6DDC2AD5C3C2052461CD9F0B7C4DECCA84297BB66C45E6A0F261FA543C5C200115A36E500362557DCEF62F31A43EA10B7D6DDD1124049E59CF7CD2839F1C0F25A4DEC917F58258F703DB3C3C096DAC7801F124F2B481B75899854C2F96A31685FEA7D827BC6693CC154AC57F2AF64ECA096575A9CFE60FB2948F739647EC82C2D53992DD36F7C40EF1A20CA46FE368C758412C6070B6B733F0198B4EAEAF192196FB26345C6E78017E4BDBAAF7DD87453EAF97819CCB4ED34E7B4E58C923FF7879B1E5040F293410DB1BDF500FC42D17C8224F0EDB3072794EC9181995657EF09D8B62B507C1DDBAF50883D7EF8C905624A3CE1D04A5262C38BB586BB2A611BEF049C4BA2EF9106967DBF2BDA2B527CD7A24094E092D2510C716AF51EB3A1DE5CC8C299A4B190A65BE7B2CF058EFA6CE01EE742A32CD1269F1824D552A45C1F72495373A43C20FF8C34BE274091229BED3787D773A3F8E9141FAB344DE560754DD4F63254E498897022C626838EFF75B4409FB8C8AF78902709FD209D5CEC28B271815763210DD803AD1EAF09856EB624E6F2F82F2E6B415E3A91FCCA0563515E6EF4F5335AA3D52C34171F15882E4B6666CB26C5547E7DDA7133F98D8CDBFC45AAA0BF8F30D9E5DE5ABE1BB1D82333B8D5FF27CF857F18206DCBA8FC8DAF0819CB0DD4D73660AAA35996174A9646CD8D42AF4C29ED82CC21214F621E80F02D72204017A250FE3507D53166A6E52E57D1EB8ABD06F94D6F4D3F31C8FDA69D3FAC67967998070F8FE7D5233C3DF64809F7FF00C68A66234391E0C5E94F6EB1AB8D3C6CE0550C1E66624BD5829E3D9BC85B429065C85CBD7C31812144C5FBDA673D57CFB5151CBBDAF7A889C79DBB4D1BA7F43C4F819E868D593EE06D1D7F3A25071F27E507B7C006F9182FF0CD3A23A27AA4DBB89567DD1F3C199286455D187E25FDC55021628E18BC0C1A88FF49A0F23A3B7FF95F48278EDBAC18462D26F63D77BBD8B5C3329CCF8C64E984B9BF960427DD794B3FF4BC11A0412B3A758B5D643BD4FE176B333FB6614715AF5FC28F0C2D70298EEACC02BE51F26822FB98500A20E7C299B8ACFBED9181CB5576DE2A8A3C0D05E64EED3227B9E93AA5AC27402B1DD7F934566C031A85E14DF7D837F5C5C31A28CFCE21AEEBC8B6D62F494A9ED5702A59D09E4B1C8ED31ADCC506DEF468BCCD5DFD774D58A367987F52363AF0A4FF151492336F66C8E63E1CD041C9E4C01AD87CA178B5790480A26780332E6AA32889F8EB853CB349EDFC6BACA5836D0528FC07363B403854BC4C32CE836C29472FCB23FAB43AFEDF28F9AEB36E5127D82556E9C5A49AC13DB026BAC273200C30FD4211A3C853B51BB7DA5527ADE4719FC7D12D3CA5EAE8595AA8F5F282058F5A8CE8B4CDF42003A5F4DE596F952D73F2B87F7A85051C578C74CB8F36FE91859D11F4F43C39CEEE140BEFB3E7CFB3BB16B234528DD4F0565E9551330B1A4CDF18BFCC3460666F6F122FD8AC148968976344CA49A4CECD0B2E212D5E3453F616D4151F85528C9A6BC352E102C2B8D1C65785AFBBCBD0A4FC05A6EB0159D071E244410125F443113B6F28A7D354CA39565B621420FA75431DC65CBCFAB5C491BB918BDD3F5FC1A1FCBCD815FF989C00258899F24C8E68A954BD09D9B3D8F1F92D22CA9B4F438A0164740CE45A8D9376C44B65AC0D596A19D9BE5C69E5C42A6010DA5B6FC95464FFE13E36392966FEAC0EB542112E394CCA7F584FF2936973C00F48386EC10E3DEB7D8C6CD993D7794971070472D9FC6CDC7732A509FFC43B61833072D3A1DED0209B71403079CF3F94166FCE366FCE702D1E7B0BA6B8852A0A9092C586D480FE53D51BA11FFFB2C54003D8D5EF2B0CA099B21B538B6760A0ECA3383744DA4036B3FCDD5C2236E84FA2D4C505690C775A7E7457B6B43BEAD781D6FB088094631071F924D585304F565295298DCAC3570A4164BF1B94393EFD01BC969AEFB7B2EB27C1A31ADE6CCDC221D39487496BE6B6A9C4754B407CF06B4C02A49E79E866FDEC53726B36684783B65E3E54F34A6FEBD96D201CD4E5229F304ABE705EA598EF5DD6CE44CEE6EAB3E34E7001B4A1AE5A0CEE741D51D4FBA32AB50490A87DF344A22A50A67240186767C81A88B567A36822B66CD1E405959B5BF5DD92E249BB52219674D7D9594E822D38CD8792662A78255FA62ADEF7F19AEE9F6A618ADBF3D13622088B1EC59BE816F8D33A0CDE071301293DE005B79A11CEB4D00D4CF2EBD1EA7B7A0525D3A08D22A1FEE65A304FA7699D039512EEEE4FB1071913415A3C40797F1C95F54705C30EC5D0044D1A3F6982557EF81C715E1DA49DC065A2BEE52732ED9596157747C4DB1C176CEFAA23B92A0F26817DABCA2CB3637AFEEF6B9BF082E5D2BF73FE4607640F52F0DC749D9E9A75DA88470D2503500A1E7E1AFA1C80F08F62EEF21FA3F02D03F3243BEEDA9202420E10C7D838162FF32D08E339014B3F7213A3BA94F8B415DC24AA72790947BDB4587E05EF26E09B8F20D19D181D85B5EC57510A50554682622185D1ED8E60D25015791350FF710D1D800D5881A7B31243C1053863538E9C82E849F7DD010B121F1014D018C79DC7C9648E115D92C9AFF76AC55470A089DCA38CD00939DEE156A7D3ABB772FFF15408AC27321D1BCF7A5C7A648DA2E51B30C75213D0C85F4D0196040BA91EA1FA1224DD727842662A2C2A720743E2077F57FE616EFCB119E58335BD7EEB975630249887896B8C9700F03D48378D3F563B8D55D163D9A92B9DB0209DF84AC05EEA5DD2C8E61DBF9FF4492F0ABEEB7AF7024DED8EC32C4C1F2A1108B01FA6C6E4DF68D1514571E9D414578228C2BD086C5061A0D8305E22D33080DF50006B64302AA87A9C1505691A69CD8D0B7D1D10FA8C0A9D2FDE265FD11D5CA80978A5C3828C29C5BF05D93CD2089B7962EBC0828B5A2FEA712533C53457A640911EE2A7AE7333BA2884D73CDBA2022C9ADD66994651A9A39793CA5B7381EF87F4ADDBB6E9A9128708D0179776C373FE005D90B7113D04ACD13C0ACF1DF2F8CDAAC11EFB8FE1AF1FE093069D2AB77B47BBC5751F50553D212306E4CD8FA3F15E93BC8794BBCB63A55D49BD890E6D96633257DC0FDB41D19E2D0919280C3BEA22AA20BFE7C1402188757C7FD3C33F38D81A8B28072E593DAF74C4B4EE96224BA3E3C3FCA450263AD7C9FDB54AFB619EEEC378958F7E0150779D405BC622A8FDEC1046273CA71742F7A2962E84BAE2AE357C8F1802E690DD9303CA83CD7C63C3B9E2641AA8704BFC060B1E8423499329980B066A77DD69E8F4A43F977AF8136A57A5C68F0AB5DDE811E1E42CF853368062D61A2590EC72BFF1CE61B408EDED1D076F9BB0A0101A7C82430BCDFB8A265E204B3BC4DD7A02D4E0DBD0D1A230C326DE75C6DF242D14E2A84871EF117731A821787653AE248773B41D9FA850450F1493E5389CBC70F0C5BDF6F5652DDA2E9CF79F0491AE7FE1C5DE3ED0A2A368511DA7DEC4C40727E083CF81978E58DC548DDE2182EC2864610D1DA7D9026DFAD28083346D9B9C195397B79678000F9237838C4CFB8135021BF03BE30CA3D8B91E0114E94521B78AABA8D892C52B67286BCD261998BE839FBC07FD04BC3314E22C18F72B19AA31CE123E59B9D8C8BD0778D00EB2FF4BD80A5D033746477397DA95570CB8F3DB93593F8DECD9EB06C9777396ABFBF8F2CA730E896A44F8A968A7456168275CA6CFEDC9EB4252E471F884DE7F15ED21A1C885426E21572CBE87E691226BC23969B51C7D37B317E9DA2678B6B84FB0DC66800F76F81FD6210586A63BA8790D21E67452FD16128477120C2437F70FEF03505D4CC63C320F498E4250784F3DEC070E5C4D859AF4BE813D96548484DA11101D41C9E325466B0811922E792751C4B2B4FCD63C60AB820E45FEFF6C0A5A63C5922045F336A41943BAE4E016618059B1BD82B16EE91C4AE2AB47FC8524B498F4171B45770DFC2C83A143DD0F1E8CBF8B0DC98F51DB14568BE566CB60DC6505E89FF1A9915DD2926E2EDF231686D6B8E82BD028B7AD5786D009A660A952780B58E79BE1AAFF67005460B314DAEC9B26F8CB4B7C6EBBF357785E711F97FB82B1F3F622F2F5F3203120E201BC18415FF86F9446B7812A2DE841C6FBC1C270A3D01C3E8A4B492C55176AAC3EA82CE2A73B12C623471E89FEC051E20438377A4BD3CAB3E2A005F2A00BD039535DCD7558E54E1259EB78FF5F94E2D526ADDC4AAF68EC6CAABE963B7C281A8C26A2ABCBCAF84F1BD7172E081E9932D58A7C332C171F272BFC15A8EFE4397FA51C4520779F301E3F1E266D96175C83EFE09AB889058AEFD3FE7906D16ED0090CD8D28D0D6F59566EB765225C8C3421D56574F11F0E51D6E95B4FC71315C68B7B4CD0C856DC80F632A76D59B4C0D5D73931F176EDEA52FDCEC892719379421D2E43F9C9D2100FE1EDD01133028ABF1FEC43B9129A2AD44BBC34B5949678B444C841B4C92F77118FE528CA6D44F8B9A1F57BFF29DD96ABFC98D726A6470E562811B809719D21B2A56EE6161EF61154F81600323176EBD8B26D023AB47D611B973138F1D27EFB4972B7AFD3B6C1418EC5D5ABC815975E69369E47C4038D4FAA13F0B640107F6C25D71AB22E0C832EEF47F1A379E536FB44EDFD75FC1D766C8AFA31C1ED642EE3B2D808CB16B56BAA4F3F198992182EBA10A3A4407F16A24E6BB047C9DA14EE2F6A7C9920B5D538C91F78DB70184A5084515B16558CF706750268DF73CBE8564E8F4B55F98700FA74898A2923710F96152779A012A589F2B9C3F38BC6BEE7854B4B57F46DED05E563F960D871E4F12BB97AE669F23C63D932697E0DCE92A54C5482D34E9D95F9F23E923ECD6FE8F8C9562BF010AC281E765B887093D19DFF0FA82CE02B82605559CBC55D7E4A060C51CD04CBC1638B0EF3C8ED7738396D354D91AE503887BB66FEF43B809C3C597A9476F91B73C5BDE44D0F06B93EE86181646CEE8AF7D6C829EE4F34AD8334DA9964B2358A29DEAE99D9B733FA63A157FD230F20E324B8E86DCDD6E3ABFA125B8F700F7847F0089856D37E7CDDE011E9C25BEBD767606D95994899F4D722289606D1791947B905CC30C9EA14026B7657E3DDEADFD49E0B45681D99A427DDC50853C5FCDCE4452A08037BA370C8E30B9C86AB2CF2CDE9B79CACF375092642FAA44509C8510BBE3F221F8DB5C5DBA97DF130F27C6D6BB017D8B7AED64D7D816A3DBB4C70A944E35105CA34051802849BD5617F32337E3A7A32528F6C118CE63EB93C1FE8E124F1AC68EE768A1187AB304B328FE99808EACC6924F178701CD5192D658853E896CA68A860827283FA2C5B8DCADF8A44785093C921ADAD5533B927EC378C773C4C667903E9003B512F15057A62A25C2C752C0EFAA003C5D8AC5B07F552DF3E85CA2BA7884D5A42A7A560A4A9978064C1BF0A28065C343F73AB1C16EA93FA06ED0844A37690DBA3B3C174B427E8D4595267A52D543A9A0B0B8F2D3ED00FA6F3083FA0D16092EDD51B54806637CED50D6D974C45DC132DBBF94DA4B3054971E1861E0411604C1765A00E5B3BCBAFD07023EBDEB07FE1B23464514848137D799E2E5E6A0433EDC62D9ACD9335DEAE26A183BEC45A750CEE5AD71FBE1D3447763684CF18DFBB64AEB42ABAC8E45399E31B27C8020921EA224C48A92E1EA64FDBBFFC56EA7A068128CEB4D73199C041FF5FAE69618586C2D9CAF8C8CEF2DB8100D69DA0E00A1C2ADF012E1FDFE12186D60057631FD925B5134EAEA66742A7062E0119F10EC518577F05CB61214CFB9473525DA14C46D4917E8BAC522C05EBA8B42F699D63F0CF64C2D172E964415BF6F21DCA8A29F62AF00B8A84197BF9A90AB81370383A70284B2C1E365382AC841949FDACC28DB6045A5BB945AA561388E625F3972705647594EEAE2200721E61F81025737D94D4ED2C9D8AD3994BEC768CA8AC7F8E5E0A3318D0237F60CC190FF7EA80A1ED8802237A38D817F992D90E138A611B431729ED9E052EB375EE53455ED26DB244BDD2EC9C9F5FCB5F5551A113FFB722CDBEF55B0B1336A1F825AA2F4D0E25D66FE5086F86F41DAD248439D585DCC99F56E2DABE22C2D9E300E3A53FC7050A620760C55EACFFD3E9E97C81255DA0E302586B0086BD4D4919DAA37BBC9F84173D3FF12F9717956DCC7A01967E4E66FBBFEA9F72463CBBA7FACB817571FB62DB4898AA02BD200684E7E3BB942082656030AA62F3111BBE1A4B83FD8AABE7D9E87B1DA284F45EA9CBF43A080556C58F2D2AF589442561C0C1E98F40C350020D0228092FA093DC8C875687277495246D155BE60D8E8600C994F7CEB33258BB37CB4F05E4B924A0CC0151B8C2F78693940C966BD977DD6ECE0B92CF3EC4B5A50D385D0F3149CC4D217349C2194BAC65B285A06B7B52D9461D963B8A712D88B93471041805575586F6007793AB34AB2E86FFCD23B532E0E4D3150CECADEA6C51A78A10AD1ACF6173FEAAAEE3E63547ADF6F645AE30B8F102EA6DA77A862D5943D9367CB2EBC5E2F73F1680931BB8309D5864C1C7B7D6530D2F80B978A1AF203CC5FBD1DA4EF4D26838B68E068CC030A87FB9E18526032D83899930AECB1C743631508FA7BDFCB98F929527A28DE9E108BB542130F4EB6884783D3578E10C4FABE2097E82E2441E3DD18FC35E17C2D4BFBE083E387C2AC91DC7D64EEA11D77A49D3DA76EED9FD7126C8F7D2883AD31B3C8F8B95DF2EDAD39FAC21953A5F7D14110B6231D4B4BA6A9B5ACB7802D9694421DCE1EBB320C44020AF26F0D62C75EB7F4CD1B73D3BFE9381FD48DA2BECB5F7E78BF4F42525403913A5EC9EB648C14711C0F3456E021D81CE4BA49F8EC58902CF65C08698530106DDB6AC65585A326EC6ABEDFA2E70F34C8E3A5F91B9E10ADCF213B27B4094581BF10673B74B69E0B68A42592B8CC8837BC9FF053E7A6C9D4BE34D3D0B6383D9B41C17A7E237525794A5107F429C552A46B6B70CABF591826D93E3DA6218BC76EB57BD050471424DDFA31B8363E9A0E0F6D994B8DA1388729C1A525E41C421C84D95556AC0D2FD89C63A89C8B9EF3469962399A3FFD79EB0E15921D0A6F011E9CC356B80043FA6E82BDC28698B8680959349FFF347399E4CCD8AB9E8EFBF7A6938BB310F4F26FCBC2E193CAA1DFD8BD69926576B5F7193C2AA269655820EB8EF9EEE51A115C363CD6A34853519D8DF405A0B4878A5DE1B1177C389375D564BA8A1A39508C1A9D500EF0609510B1D0CBE635781A07687F5ED42E31B5E11F0553AAAB6CE586D014279C561268ECFBAD1EAFC08247397498AFA87A55960478AEC3E70E68FB87955D9E765199B83C1FE3924B1902C5A409AA79FDD585F27E17193F9CBAB7B074B9858EEAA394DC58131E405467521E6F65CB7BF35D0EFFEDEB5DDFA1BA5717824F1ADDCCA584D7A407DA6D967A3AA5A33CA005F2B9BA2D85772A94189B892B34C471BA7D4620BA9AEC7DB2C5CB28109B9F79173E5A19F4411E81A988E1EC5604C80B9C89ED17BF28DFA18686E9603B8B88CBC7849057E62B3E2264FB6CB9630646E42A3E59F5020B4668581D2982AB829095737F006F32925FD9981912F4B11B34C74A42F857A8AC177CC12B4898B3C65594A557A99FA1C5797D86DB172ACB1A9C982F8E3092E4BEDA3A4DCA7120791EC3C1EC163DBB93A4FD3775E24B943E76B387D386DC40E6517A19FF8FB6EF0744D48631CED5AF29412B91FB51D2E2D96598AB6B43CF9B832341DD1FFD7C18B0E3435C7CF966FD6C4FF5F13F8E1D684B9E81A7C3A5F766CBB35DE00C225323B17CA9A32507E5A9ED2EC34713702D5FBE5D029E748389715BF1E9F294CD08EADB2EA1859F887A462678A08FF8CFED3CF36183AC54040FEAAA9E3232452834CCFB8DF25967D6FD7E108B64E46D8E9C91EBBBA46FF53A8E1C6A1024FF30BAF0485E975C4FA28A94F16ECD9A0CDD7EB3C8977267767734CAA33C348015E25E84FA801093FDFC3D12E96B6BE9BA88DE54269F0D3D401CC75D167BC57000699561255919280D9A876C7E1FCD067EFB63AA5D8E5EB1135E837AD327A2F7DB2B3ADE67DE4C131199521FFCF061DBAA042218831F19FEB415C7D2E1DC423974342F7349FC292E46725AADB81FDBF932D7FC4297DE18E1B70103530B08695ED79FDB6A7BE8E0C652902C30B9C174EE7925BF904E5C5F43B7F1A96894EBB48C3CD465E173BFD094D8376B4CE39359E6878DD04D0E5516A8B5E485AD14909C680222A7092E73C4B835AEA5E0B1BC9F463B236BC3A5B47243F032E9CCDA15137CE735E36BF32BB8A58E1D5074A555FA99C824466CB98FD06083D42F4B43CCFC89FEDABC16BA28E3A19AF1A4E8A26A22C245A7D04EF295B5B0EF41455FBFE726A4234E5396552B504751EE74BBE14C500350C1789E99931B6DF0279B77575E7CF31BFEE83D02B922970BE3C8C3B3165DF42C2AD181B3D21A7435B3FB30810EBE90576052404E1501F6D933E9C7DAA1A51BDCBB7391780A693C1E0023DD1D608B639BD54DA8B270EEF35D001DD61305070DC8F9FE16FEFB1C17B60C83EBBD8AAA4110C33D2FF18D29030F203007DB57138819F064F4F628CDF1F4656E133C319954B8EAABD5C89C6C24183081AA1A0962C4DDF759734CAD3C9194691E21B94D5AAF1275142195171E22293393D3B3D3C7112060F8891236BA6BC3157247E3175C4CED9A7DA356AFFC5C00607E6009A5DF444E554A34353AD3D65D7C12D470B13165E473411EFD9C6D3E3B3378B534F9052AAD2BD424A0F8776FAF38E68F02357B0FE590FF54227A4442A18F264CC0AB74D30C1E6A2B736E1E1FA8CC23748441624A68FCBE195988F0BEDFB5C306952F0B3A45C8B78BD0E6FD1E874C11C8A87E3DB4A097DA46CC5A67A81CB0DF9AACABAA5AF5694B74A4272CF6041532AC3A01A369FA585116CF8F203C25FF0745151AD129FDF1338D264CA08139698341350F6A02EAB070799A316CE358CFD44E0120735C368DAD616F9B6D1251A20B40D3D3A14255C73E5DE0C2FFF5C26015F2B9A9547F6A95259C60C0AD4D5A693349A35E5E27C1082368A7B5BA0D2E58B58C07D3C630269AB45372857ED601B87CFF5F77AA0D1608ADE00D16619BD55895593901232290554ECF7F3BA98F30400F1D441C74CCF0794635AA1A65F0678E5605DD1E260F3A0C076B74396A92F798BA1A1B24793E5FAC8925ADD6F5FA9DC92FD54D8058DA12E79C9143E876A54BE54E32A5A0BFD3CEFE7356D8CE10BD4EE88082072C9E9EF3D8A8B08683C2A8E1103FB90C8F2FA9DA58C7696BC3D272F83DA7A76F18C81B1CF415F282AB2B47CA4B5AFA067DE561B9C72E86EC41266E0DE4D568A0800AA932B7600EC07425E7C26CDD3F637AC29AB356C18CBAC6769287468D281388698166441751E9A6B4BC3D9F76764A0281C18EF966BC4668982A65353C4AAAA44DF59E81E50B22A6FCFEAAC4A5368C1AD79FF2A9B4972DA83BEDD33DF59A6C594F63807A3A4892C804FCA85B9EC4C296B2FF20239494C6EA9140710FBBC072E787B36D07476D575B35BB7B4122392C5949F10B384025E7825F1EA395C2BBE998351F2104EF1E065A08C714B782FE751110097639EFD159C8F24D6D9713BF2726F3972802C707C29F160D6B769AD1D92DF1957CF49EA0CC5357B3528F38A634DB7A7C8E6A1CE5DA5EDA4F260C7DA9C84A04F94894A309E274B76AC5E2C5553E9ADACB817D3E7E2A762686B047993C7ECF019A8C531D2463B6FB2AD88EE69C838A98CC0FBDBBEB05A4CBCF853503DCCD2A89B7C4A8EAD6D0C52DEF7607C03997D0D399F2F572CDC47466A85587B65FC41B47553C9A14A7DBA10DD4641B07259B603D812DA3DE9DC300DD6FE151035A7B9024E793FFB0E53666387D2ABCECDF0F75D991EB826206EC070F2A575CC8A2CD329B2712FCEC6C5BED86B1AFFAB39957812EE9CAD12B1317F5E50FB8D0E0B5124D6556D7D3474069C0A38A68D78F33095A8C662B85A7D4C15DF6200F6586E15C9CA5BFF33C5B4764A71E4C96CF998B42DD51055350E626CE38AEC83F906EA699102BA74F1419B5AC3D96E53652104C5D502BF5AF6D08A83680E8E3879CDB25E6943B6950DF959F4F2EB9C11F15DFA30B112950E48C5CD791E89AB90FEA28788E62231DBFF9D197BA9A540C397E3B5DEBAF2F948ACE56AE6D6A0E8DE5BE48C924E6089EF34FAAE96D1AB5531843804544C211D835514A63E398AEB186119F47A051E3AB8CF89CC51234E6E985D464AAE3D39BA96775B0FC9B06396485407E0603EF178FEC94153892ADABEDDA50D1CFBE3C65C87E437E4998C05DF4D5659D80B81A257B731075A266CD11F33849ED6CBB601EBEA2D79BCE39F73E2BA925CDC6AEF92345D477F545975713FAC7F5CB49A036F4818215CC10E6FCFFD437F16C40E89F87C7D7AEDB74EB24CA317EB15C78C8B6DD029982C1B772EED57ED81A2E6A2E7882202F51ED3EA17DEE631D567884F3607921F3936EFE8897C610F6FDCF8F91655B93ECF6A2F1A61EAC4E527AC20D142ECA7644E6E90045C085C7AD3AE96E1C5D501E24A16C759BB0A92A84EB2DDA17AF3DA6057E187C86E6B1B50E9FCE71D5B5D7AB9F0E7A9B45BFB3BFA47518B78253FA35228912412D4FE85BEEBE5B993EEDB640FB4A7B0BBB956FA45764748F79C9D1898D3BE690FEF84AB66A2FFE3DE7282608594ED89DDDC9278B32336B9C538A90CE0A295164CEE8B602496A0D1801C0F74B5C9D7E50E3E842466194ACCE6B23D7D20F914F13B1134CD49607933512E029AB077454F8A7D26C007116C53591C2295DADC408665511344987DA2EB549BC3B9976E20CB4B231C8AA274925119E492445F8CCB081BAFC532D5A17F6F8AD579C5E8AF825BC5CF035D830838E5522A0A89F5B7FB4116F80A90B33553B6799C6964CD271E976FBAA84A18B9D7E9CD0ECE9D94C7DDECC0FEEAE550387B26A83312D6E216002A0F0BCE93D7A421ABBE0A371F21A41BD4D295C6500649A7EF055F164A4218E9FC6909C6ABC26558EB41F7A87BEE5F426A1218461716768E610D5EAFAC2F5596F0DA32056889BEA04E756381B5EA4D41BFC0D0DF96A15B8CED05CE719D1C44717985E61013F1920D43B40CC9F1646A63829BEE1D61AF7CE8F3C4241824FA7475F7049D62616EF5FDECA598CA651C3FE62F2077F48A5FD2ADB81316CBE0597328BA11CBA46CB83CC8A2001FBC6BF9348C948D55F91D21E5C5677DDC0D652FE470CC34131F1D74DFDF1165E85B1CF3EDC0D6B016877CD0004AED251371B7FDABC0A6C65AB53B4D86E28C678CC9F9E683159B6A35C25ED963526B099B429D7808AAE263D78AC734B917B8B58F19D01E6A6E8A1B9AD8DF966AF74844C3D8545EF0324F0B72C617A5036CFA6B330CD350C9589B5C84AF86A8ABBD52351E82C2E6874F3BD435A0FCDFEF8D00EE3B664E5CB7E75E3F71853AADE381A5DE89817F36AEED5A61BB0421B5D747E6D3A2531061045E1641579026D869E19BF6C3B5E01C96C6EF53FAB39F415519980CE7A88F653B00929EFB8EFD6D69BFAFE85E9A477D5650C6795C3C1DBB183F29436D5AF3E910C3B3B35ED54D951A61EC7E7846C168ADADD01743CFCABA8C51272A647E2078C1EEF2A326BCABA3D680339F430D3AE9887CA5A7B5C6D22814705E4802184CBCE3B99C4E8660E2A701459798195E67BBB273F35B661F1A245CB04C302AA49D3DB0B6DC4149E674B6351D90C6BA9F6C138567D2B927155E7068944A73B7B98E3FCB91DA80F20B32AD6381E014EF624B97D7C607C0C035B74F7427E6091ABC885C5B351B19179CE58E2D295DBDCBA3A7A5ABCE4101B9062E18B77D9AE11E61F59668DADB31295D6E8014910CE63223FB36C4F7D194ABD2C44BE6D0247EAD4E8697E865C563D0736EE96B0EED88CE36315E13EFDE5C48F15D84F9A0411C86AD962BB8381533034CC46546C8176970A8E3E2D5FB03A444ACB317EC9004C1A5039CA6BC2EE2E3FC111FD4E6610E006E66A047C31E795F75ED1008A84771C77CA73A7D88A5C501498CC4BBE49FF3B09E359A4BC39B67AA7550908B47920F78010284C16003A82CCED9FBB3F8A1CB66F88D843BE4C1871E286F02A22A7040F156BEACC4854168E9E9A8BA9D1FEB474477B55A82DBBB5ABEE97335E5FBF8190061700FE4BCB7D9F1EC643C39A4754B63020EEDAAEF521E466DC9FDD1146DB60DF51621A0FA11BD9C8F0166A805067EFC4D975A1C0BCA8DF5C5A14D2B435264D2881C18294EB254966D0CD5840CCE5050EF7FB03A48670A265C3C086DEB09EB4AAC34D86493982817F73382258F613A53A741DACBA1774BACCC9B2C89F3EBFD71984DFE4D0A6F539AFBCF13BC830B1D4613E9809B18A4D1663F56CB9195FE6776F503D98165F910F8675D013F0E3446985EBB1719F8CE920CC6D9FE76A881B8D9433A9004FAF84E0A2B41164DA37C5C377B2A3BE314C7B8A74EA8384E95F9CD4DF15C11C1D0A5A21D31EABD6989D90FB327431F848FB5210369EC8C76F00527247FABAFE9DDBF9FF830C733B25625E31DC415971D33954FD3E0A094B486223C83518A5F39185DCEDA39F3176CEB6E8B12C4C6D38F476E5542120F85AE8538C9040564563F7CF650BBD48244916CF4B6A023F3AE5D54FBBD94CAA67D8410021F6613A7DEB9D823DA04EC92ABA3B3DF429BBB5EC0EA79653CB629DE8F2951ABFF2DA611217A8EDBD6B1D1CEC419FCA8807CFB54DC47797C8F39ECF834346A8CF56D49942880E8E81B4542B2675517488F620D124D5BE2B82794609FDED401E7B2201667F6A5B03BF8F34FF90491D25CBF6C719D7105E4633BDFC3D5B346191106AE79779777801976064870984E28D08C593C9FBA45E7E4D538D29B9B89CBC9228D09396A37CA87542314ADC06579248E41A38C698EE5A6A42AE8F1A4F734C0083917EDDED34E965D3920A65F44A099AE2E8CC10C051D21F7877DA2F2723106A4B4B0201DFF275CB0B5337DA286A863949C330A826F23DBCFEF533BE979AD5249554765DD65824FF7AA827D3B9EB27E326CAF45D80419F88D69891D568DA3B0C7469EEF9B507E59AE5D227BC32CE9A60667174FB4441952472A0439C406F002224BE386E0B6A6C73699726C333DAC412A01219C95ECF601EA3DC5B494436724F1EDC240C221C9F76D6522689FFFA455365D6A1F76A64D85C12BC5412DB3F6E178E7E2BA6E521D74715EEB2D6E6A90BDFC689E6C9FCF15503F647393E4F001D986E3380497EA85A1227A6E479DFC5672C731F2F38400FA0970C4EBC9DBFAC0AE5FA891E7EC78AEA8D26E6C0AE486F163AE6EFE829C3BF78F9AC3A7233520012A85DA34B0AA617A4D3398345EDB3EA9624D970F7E0A153A63EE279CE5B17536E7F93582FDCD282DD22E2EB25A5AB6474591495F3AA5AC835DA6CECDEF125322428B4EFEF139FBA6998043F94FC5A986534866B515CABA452ED90B25BE132CFCA107A66A63A3D2C9AA8DDCD8D702D9B3C1B05B9755E49B95AB8DBFC1556E4F8979DCA67E57A02798F1B6D53D88FDA6976D040BE1EE6D8F59A596C26DDC9F912BC1FE74A712C30D3B9C94A2F8B0E7CB614872D0742BEB599FA74F7D4D11A095508F4CC0280F7CAFF2B3F9C674E5A08BAEB4690568D4D57B6F20CAE55521311FBC28BAE3B47A5085C128C0F04C50ED04E2F5609CFC04B8CCC7D2DFF776986EDBBA456BF6E50B37CF252E715CA849746C2C247C8675E836E915C5886149CE5D8687ACD21FA239694128CD0CB380739AB41DE66C78F6C1CBB3E15C61B6BF1C4EC97D9CAB128B32943574DE1CE4F4B867F78814EF4039681655CAB249F671BFD709FF3F58208862C8B8B9066730C09E9BCF8D6D5D420EEF2F414F16DC5D3EEFD104F0AFE8718441FF9F1AECD96E4C76967337C8590EE8DE865D970CE971A0555ABF92A1F559BB260979BE950FBF5B55534CDA139B751D4A74A292BF6DD8BC4E183E8C16A78681A131D651CFD8742DFCA60B3BAF40AB4057E623A449F0801BBF7D63B67DED5B4B0B099FA8A48CBD86B87392E85437036DD2B8A4FC27512A3DA41BE300B1C332BF4692B2059686FDCE04DF947C9D30D215F08420FE9EA99A84CB98F09E30D03EE3B8EAF63AD60F6090C7DCE52BC4DC91B5FC6E599C24E7EF411BC7B989E3248554049B608590BDBFD9A72958C8010A734045C2E900548546A0D80A93543146CDAAA6F79427DDA999ECBAB120783CCD57D1D481407E5138F05DB2DC7CF1E964D62501F0C611DD338677EB3BC32EFE2AE10DDF3EF1A2CEFE71753C2AD9140B56D13D07D3B8DE6D2794A50F7BCC94CD66C2DEFCB2F622E509E7C63AACAA01449DD2E57B085C0C8CEE8E3D304D2EBB61BB46E6F2A69A3C2011C4C48B821EBB2B24BDB9650E4502F40EE3D7B2E03571280E0C9C441E5B2371F6561A300A7D34F839DD01830357CEBBC6DD6002A02325EE645183F541CE179377F472B807700E69498437836D0C1A8CA47F8057138965D45ACD4DFA07694A0862100BC89F2D3DCFB1CEC66F9A2F57CBAAD7F9C47D6CE30CD83B136E7176BB50596EBE60A90D016D35D2AE5205356DEE559F1258B78F039D3B2B9D57551DFEDD545D16D22823B41FC557212884FFC3F20C0459CF56B4A6DDC528985E94CA5AAEF7FB7F6A866F9B4BFDC852C86A9B4C5892D4BAE8FB37307712DBA6AD622CBEC3D9CD7C40A9077E94A12D577D4B6CD3884EBAD5E171D5C58B7CE29973CCBB78F45047405C2F39355EA96E8C5C53C27C4604EF0B0C86229364EBC15CA3FAFC93A58E59DA9C816EA384DFFDCF60FCE232AD8B313E6C7479F34ED09BB95F8AF2FAEC5D7F305E8E8F97859C695C80C1BAA67A4D7B69ECDD9C1F9A74733D874E55C8730AEFEA76DFDB0335C420AB9C3F113EC8899B28029B43803EF152705D7A29E75D60EF9383B09FCBDE71BCF549124BE87B9A59F74F3EC45AC8268D771BF4E0DCA3369999BEED82985B2DCCDF5912288F964220F8B3C8ECCBBF123F9F460A25DB66B22A58F3EE6FC050AB460F5A68128CD0919724F326D27193C8B85DB16360B50CF187330B1A8E98459F7879057D76249EED2F400E0D68ACE8357695800B95861A491F7543D690F745268AC228CF752BC681BB1218573D976291A69B9707970105589995DEDCA32B34086F56BC30CB4780AF986D485AFB8C888E0BC688BB44B4EBAF0CF1C45586A65ED7314A4E295A8C848D836B1AB75AC1B27FE8605EFCEE1543EA9605AB417E22094AD4170EC65B5AE079D6F3F145B8D564D466EA6260C1CD3E2D25D3EAF6ABB97AC40B554690708E918E7FA5B5159D7C1D279E5040D9F498677AB01F8D4532085DEFC756613A4910CF2E30EBFCE8004DBB13AA1AFDCC847020B47F2CF5A2B32A653FA6C2FF600A0B6A89C93E569C1A955A450D3F245F49529D05BCA6BFA6ED6EB57C87223286A8D6E88886998B3CC15EECE9DBDC7B1BDF6898F3D4032CB25495926149FD4E279562928327C924DC7D39ECB1820538F168801F26B19DE31147DF6DCAFE510D608A1B787B7F01A420E6A3D4DFDA8A3C55CE1A3F0FE2B0322E3F36B8DF4A753BC0CA4FF277E0F906802A948C4DB5F53DAAE000C98D4E1254FEF305C2A849B68CF569DF814182379C9EDEB053883B918859F56ADDD63F68A4284C5C2C68A58CE14C4987D3549D766E03CB31BDA3A0BF172880A8B153EB62060EE3A3EEF549AD933C2BCB4A0BDE678DCDE569586E5DF98D3C1395360F1114A8AEF1EEE992C82A7375B6143293574D9D7094B12881E230F067A506D15E10EFDD186AEF6A07B6FA69CAE716E3C7F08F62D26B0A6DC4EED257F2D1A2D6999D36042730F8274114958B232A4D2A6EE528617196B39EDF2CF1C4939023E226CC1E1804DA6E39A7DB22510FA94F364E1BAE2154B384344839389618397ACCA0F3CB626CDC48D00BBBF81E26DFB3CFEB49E01C684C428B8E878E38C98BE42CEF4128DA8A920976DC16720C34A29B850269EFE66ED24A23E98FB7BB3891C39023B86F34CF1A2ABE32A5AEE6F957739727EA42DDE5B723DA033FEC47481C210A25CB28D4819ACE326074741BF9E2FA3AAC49CDFB2706C9385A3B3BE5D7CF84F24A578AE98F23BA20BD79A85D10BCFEAA37D508D5BF3F8BF8CC841C72D08A28667BA066A693032516B255EA464849D1AF81D4CDCBB86C2081BBA4B09E6A0567EDBE3D7D95F128CFD4C43EF79AA6F597BD9857295F5D28A72ED4D2EAFA4C372ABD3EFDAE62D4860AFA7D11E7903E330EC647DEC7441EFBAE9AC9DB8195FB372599F99730F089AA1F530462F38457ECD025151D704D59EB10DC3781C347E21088685AAE1C5F6C72F7D27FD9D38E7F8277E9E07C075587D8686EFDE8A4647EDFFEAE29B0512355A18BC3499B3A67ECE03A9D2154D98121CB9BF2A5FAD7B32C77CF3D9A855882ED2D8837A5E7A420335223EF325833D052B1CB90D579FD8ED6715611F2177AB74ACE2C5D936C6B6AEC046D248DF7EB0A24CE0804489F30C4418AC1932BDBAC93D45380B1546FECB9D6D1E7277EFF13E8CB8E580719AA164176E806F20D277C2E0D77BF3D1D2807744527933D0710828B909A9DB95193E46084EB478BF6EC6CC8CAAFAE231286A29443E90C389ABB40B0AB90C7CDFA2972B2DF60FC5EB4B39A3950683613D87AC49E8DBC3408A99C0DAFFE7A8048D0C33EB69EF45016971F4AE39EBD470033B76F791513CEFF94C8200CE683CBB273A8456A13857A83D19D1FDACF84C48DCDC78D0DAE92017F8107FF2A4C6EE3D909CD0396EEC920996273BEBE5D1678E5A703F41A8C52A56D30AC9B035DC917034937659E284CA3812F3B2F269999F7D2FD0ED70C2D9A3A5C2E33930FE60C2E5DDBBEC8A5660BD882802DC077838BCF243154EF1D62D6E4F60230312C3F154FDA4CA4D10422649CE9D8DD92A29F5DC9BB5ABF5E6068F6B43520C0FCF1C817DD88A9982110F3ABF99AE93187598C516D854017B600DB3ECA4339F6CBD64CA835FAAE114B372D35F146549A3A8FD0537F619017223093627E6E2056092E7F72D8B23DB87529D93348AA44B0E118A6C538E867F357E6B9CD50D559E60400D477335DFA54304327EF65FC91F8949A6E5F6809316D6C0CB176C93573473A527E1288A3F486613DE349DC2499628035F8312F234B83DBA3B61850A227D4F77AAFB2C3C988851179635262DA13D4E026EE092E4B06E16BC8700ABBB71E9B9264CC0B0B326AF9D4E8B37CF3D9DE3AD3831D617CABD9C34C26C2196C85363FAD51041476970E13D75B55478B8CD1DF3DB8CB0AF074B15CF4DA56F91C1EF06D73F583810324480F328B200EA5C24B87A73670888C16D5C0E8DA20057517FB7F785658580D5F670CF12778A801B58B41E97D64B75487F9D6575F65B1AD45A2E32D4ACD3DE758D8E2FC7A322193160D49A2C7312752E168E49323EC821686F2EF2F4C25ADDEC7E74F5FD4BFC6F25CFAD97D93DD8A4F2BE69ABF3FDF9F9A682ACE4756F7B952394BFB8D54702E60E2858F01EC729E5498B69E57733B9851FEFFAD69D716749D3BBF8DAFF7FDA05EE1D803EEAFAC382BC7D2C76B060CF0A7BCD9CB111B23BB28E60FBF1751B134CA052A6562CED50CC68337E145329A13F84AB786848E5A50DADE9FB661752A55E31A538C4F0A3E7DCBBCB72BBCD9F19ACB40D7D226CC6C7057F33121E266F7A0E82A73C3508BCA61F399D87C11A2C15A307D30F418FBD595D8AC66E36AFE9BC4FE4291C1EE21DA7EB5F39F55094BC55E732AF16A958E2E727AD891809BD7C3E265976B6EC0824F10AED5569A570E8E18E83515B80D9CB38FC8F29B73CC041CDB1862A49ECB04723395496048751DE97C28FFCC962B5C9FA1CD082D1023EFC23A675DF1768ED2B8A069CDCF164CF94AACA8E2A9AD06E0381FE962DC2B2EFB4A5238F5277D8478F653CD96AA4AA2AA212C40FAB2325D1192E525C317185076BFF001759DC7E3BE1F3AAF26F3EA9C3F154F1033A8273D6AB5089D982A7906991BEF20616B8C785C260A85AB9DBC5285670BEF1797667828142539BEAA7407F0CE965327FFB9912E581E077A55717C626D01DFA5CA3E338D84F18A7C93E42925C12D2B01558122FBE0071A283F2986515424E06B11D9730D4E5FA431B081DFC8277B557830EE0A16D6C355F11D5892184A36D8948623482EED9EB7B70A2FD2513ED429B5CBF7631618195DCAEA035063B0D0653F805584C593BF5684B0507E8625722CA3A54810EF50C433161DF2C92D5549766DAE5DD68FB93DE73393C73186C045E5320CFF4D63F269A20F7D504916416B9BA4480CDC216911E2490C7E1F2105399014EFD0B4F2D83D8EABAB15AC4662358D16B56F379C2347D7BCFE6F7C2F8D48150B006C7AC8B8573D8E2709CA1394756126EEF317555A3D81BAE1A4219CE0FF97C42E7C42CFEEE27F7BF00CF9BC31359AF74EEDA36A1B332A6A50A2C3F448006EA79A23A9A115F4F7E4DF6C3AE0D6E491CD8B314F26036E24E56B04C5910613403B070D279E5F1A56DD9D5B3A8B493C423792B595B5C4B5561D1AD574B6C7C001BE617435AA51489C6738B4B33FEA5E3212D989ED4C538735620550EEA5CD91EBCE3A2D5F5372A0D217A6031D99CE3598ABD98D017995F623C3DA6D416604CBFD162C6AFE07C12B0AEDA86EF002393CE7E0D394933B50E2F8F262BF9EF03839AC8C53D9452FEC087658ADD1D6F1C523E98A386F1FB2F56D6C1942701E0863AF9AD5458846808259411161DB7D8A77404412B51D8813572BE4D828BD5FC116AADC5A170916658FC49DEC61C5D17AE9C71E54C440FD6CEF8C8F632A529C29E7B5E5664FB12CBAF4A42766B035BE69CC8E1A16855B7A71FF4CFFDB3140563EC30A98C833FE1E6AF596E9AC80AC3C44956A26EF4971F5FF35E153DEA3C94D9B102780AD5C17722748631A5CF43642BCE3D2F665959B2430806B90476B5C09D4862818A1086D8341AC7903C72BA427D17E0D335CE8E4899462A827932161456FF5D1A6382B86078CB9592936C62033A443D074215A77822E1ED003CB1D6B51B0B17DA10AD74B3C9F24FBD8C579315D6EA7FE46884E6C51578BE81F01CF64FBA48FC8B98BE653FEDE1975B22742FC1E418A6D1DD4F14733971E5DAB3B3209DD5E41DDBBC2413C99F7B0481D13DF35433CC13932BEA211B8F4F8B7D385AEE553E13227CCAECF4609599C0E9A724DEE75E9AA0B209869381AD40B69ED7A4F8C7D7E28849DC464685EDBBE297ED6555689A50A6223D18EE99B77C1752BAB2B983366549521F83591CAEA8D11E1C5F924EF0E4115D9A3F5C9EF3D3CA9C8F79C1B891E04E1E5D1D54621F9C5F3C28365A8DD97B013DCEFF2D89ED3513AD121738BED3DE3AF9E384554CF8E7F932161DCC295E5E59BEFB50BEB7F1FE78FFEC7B933D45DE5CDDE52E0B7C6C8872A1A28FD8A956E0081060A1BDD73526FBF5C6082702A3D51B9337C09991148EE860871332A7DD597E278F3A62D7980D464D3D164ABA7BEADF019C07B2137888488F77F5DDD9BA9C4D050885BF1A3CD54AEEDD8C4E174049775F88712AEC3371E35B7CBB32C6E01AE37E328ACE467C7D2AB82805B66E88BF02B776777A9020EF1D2B5DB5EA2C660CC594C6FCB85705DC2126817FD599FE22CC9614820B984C88B24B92053EA84DDF5B4416896EAB35135CC5CBBF61D15F2A1B5DAF6B24D32B2E908DEFFB84E614C8E18AD8BFB5CB1B72DF14A9E47F5DFF170CBC4D229839828FA4AAA251525CADF2447D7A89E4DAFFB80491DDB96C6E12E603EEAA18377F3A0D5AA8B33DE1AF6DAD0E268793CEE58FE050BA12478FD1990D23E8B4C58D2B88E8EC12A1CFC82406'
		},
		SiggenCaseItem{
			tcid:      3
			deferred:  false
			sk:        '5220590D3EFBEDC5695CD224320FDC910EED2497A72AF1561B35169BEE722C055598BF4373B73674755331C6C06225786647598C28F11D41F8576EC69913647F'
			pk:        '5598BF4373B73674755331C6C06225786647598C28F11D41F8576EC69913647F'
			message:   'D946A88701381E810269BC9943289A601521407E7DD77D3FA6B87018645395EA380443936A1CEF9D44035BAE99CC01EB6A15DEB45651651DDA12A3F0D562855E18556545130576F3D697D0E2F558524AA9467BE9B1AD409E4A5798E110C53414E55107EC17AA31E5FF8F6296F0AF7473F4B3B60A766BB01F427DEF44EB7683382DC0926ACB46FE5F51F15562CC821B399B835793FE62D577BBD232160A82D754F22F180BE910F64B47B46D4CE36CF17493F9C7C2CB756746CC7B7BC2914513BE3D38CEBEF6AF336346220865A8A1F33794C45C1D41158DC0ED0FBB1C743D6D4F1915EDD6A38639EF1708D8583555558798EFFFFF952DD32B0E7145309E4B6C1E7A3EBBFE298B2693C4F14B14419B32333F5A68E05BE88DD5131761C91AFDE1631D19F4688895E100D05AE82302E742703B5F2E80AE8A386EA643930A8BF6EEAD154EFC840B6D926DDA166B93573418A721EDC009ABF6B1199EFFD51B03BC163BEE40571B8E645DFC68D97760A4D66E7C5E96C6A232DDED6C698AE9686AFB4752770F6AC6B0773DE88FF3E799631BA4876840164A0E8E4A58060793CC4DECEF5072DB7C495DD7BC75E1D5307D36F474FC573655594BB92DF358C79D6CED1EBDBF701D8DD818FBBDBE9962043B81A320A47480EA0AAC606D00B395441B9556D8E510B2205699E97D414101B9B9B9E0889DE233C2C504CE71917427C1963DFFBF531CBE1C0A4003D83746EED91EF1E227742B821A55A9F4A32CBC615A7120C3301A1FAB9BE155B420FC896CBAA7FB2EF2CE99E2596E19DFFEB79F71BE600061A30096D44CE4B0C05785F13335A8AC439E7BC25AD3C4C4C7EF6C8F4CA2AC391130BE1466EA99AAB4286CA61E35084B8E04411EF8713020B867816EF699D92DFDA3263C8136B084BD74338AF47C2B485D622825CFAADD376D3F4A166F561EE8B36122497E66AEB72911C8D6A99D60037DF1C515828C8E20EDA4A230EDD996854ADD28547FA9392278ABB25ECACADC0F6F38F005DC69C6DBB5A2F3B7882762DC6F93A086ADCF3B6EF7A17E486843C3E05C2B5750B60519EB63D624BB1730C4F6F31BA28DAA393BC789A60BF55429B2D95E0BE84D1E55F711214BBFE896C5150297D2711A1D21EB457875A6AD173A3622BFBB802D335BC96535BFAF967EB33C2F5423308A4C7194DE381CA8E7BA2DD1D0E13E9CD3F46925C75DBE8BB2FF2361215C60DAE90A18605B8E749759232623C172AEBAE0D599902E0C3BA3ADCC2353CF75CC0EDEEE437F9C1E716C84983102006B58D553F3D6ED6B3EC92C8AB47FCDFAF92F8A26278E1A4702ADB7C204CFF838C5572C991D4CFF00F2356C088A8149D6347053906AC85898F2F3A0F2D7DFA1ABD1B70CFE55016B4CC0F5EE80260C3AA2A08EA2A57AC9F0D156829B8999BFF5E0B59215C524E964D616CE5A5A9AAF1A8D7D39B2CDC0573EE77D30E8BAD7821A1A50882F419AB7DC525B62FCB8B06D023E3D730CB4DA4669E5D4AF7D013CC03913860BC89DEE580089EE8C13293C1296FA31247B1196A12618251D999B40CADE6E8C39CB47673463B884A255005E8F026D4BBECB1B2FC54C525330D15111852B448D72B93E7FE2B8FD3FABD6E3F37949F76EAA206C0E6CE145774B292032A3645B85497AA88670176B2ADA87100BC49D7D5104F475E0B18D071A3FAF974DE3D8C6BCE2A791F69AFB631F001D9C74FB8527E277040A69203D2DDB714282D3376C4877FB0B91EB80F4550F5E951EDE69795CC283CFBA2C4FC2C7749311EBEF0AC1B51EFC05ED5748AAB232305A2CE8B1C0EC5D328D95ED8B457DE963D996322786698A7DCF9F55D68E5018BC4672CCAB2B4D29431376744C33EE9C5BC4E598C26E78A327D713FFEA2F70A801E1207AE1D8AD497258A09F29906291CF8A84473652F9DCC053A55974C082E3B29F05AEC4BE26E00B1CEABC4B38F6CC3187BF6C1323480790E43908B8B8655C15EBD8205D93188FF7986A7E598AC1F95C5D11D91C97CF8BC06242DD4E1D78759B43460C32522A4261DC04E2AE0869D2C18726302E00A05CF80A7387D67A6CFC7B1887C25C8381828E40DABCF4C79633E91857BA19F38E2206A38FB3D4B8833B99F9AA443B53EB18413F24BC22A6FF88BE48405AB505F5255DC216479BC2C1B2FDFD63F350547B2A720DBF0F19EBE41CEA2B76966B8038FCEDFA99B77D5D25014F3DA807C2EAB334DEABDBEE02E220F67993A5C1C411F0A60426DE03895AD54DFBC2F23AE25EB090ED3AA85B273D22CBFE221153AB21C341778B66737AA16F8707022C25AE1F198BE651E3885268316A9958A5F8E1DC5028E7A059FCE997E1D0C2FBC458A8BC23A31BF32FFB4AAAE1D187500A5B723282CB5BD5E1D1C3357E164D2D323439B8BBA3B3172B63A8ABFDC8721C3168AD2EFEF52FFD11635FD7BA4657D7A7477354EDB8B8B8897027B2C86C3840A97E7CD5EEF475A6892771735C3D875216701836091B9AAD3E9C22739BB92483D7BB1542996D48BF7E7C708866F654ACE4C36BEDF010FCBEC0154237B3F322F9B0D76AB1E96B16815E084705DA5BC381D3D567BDB2D45B426CFEAEAFEEA7C7C5824AE4297728824B811DC24B5269BD6EC531DE7AB9A4439401E2D96BB7979F2153996F97CA89B2B2502062F5695C24466A65478EC81B5FF1E1AEB22ADBD26BE3132BA876B028D40DC0A69618962442B40CB53E237BB24CFC101FBF9E967259E638F81AAB1131FCA988C24014186F11A14C489D34B9A4DC2DD7B9A8ACD15CD000BBAE88A7C68EFDAAE9F7C757E023B6B8CC91FB66731494C0A0E03A0EDBE5A0501A2138CE28DE3247AF11484D657C0E11C8839272ADEA22F47CB086F8D6ACBB32452DD4EF357E3C5E03A8509608117126D911BB9718E67DEE106D4D643D35F000A7515FD6A3E722831BAA582AD93361CA15C32EC7AC6384A40377D6570257095CD32AC96ADB86E907D867FB9C8A8166E7C54FBC4692C42A71BC3A5D8DEEFBEB1647E3AC3F1A271AD20AC08BD7D540DE6104C553ED6E513F7F69E391F558F4C7643FD0DC69E26BAC183D2A98D14494554D30B681B6602AE7244C8EAAC73F57FCA291D06B2A8D0F17867CB31855758B0E14ABD14D55965934AAFA6A78FAF128CC557F0D5D52A8001E7D0C181095D4E18FC5899CF00BAD7CAFEF22142AAC8C239E8C48EC36045197B19BDCFBD2464857BE2517051E90B51442B611AEEA5A9BFB79DE5E58ED9306A6CAA72DA520F033C19D0D6EC5A80502FDE535803DAA1B3FDE40FDEB0508E6652DEABF0B208E9A4AC3F4BCCA2939DBF964E4673F52C0F165D5C7BB3F6BB3287E6836A8A1A16AE6652487412F10F1069A7F689F2D874E9BD58C607506F3BFD20424CDBB30D45B610411EE8EED967EC64BCEAFFE3DB84C4C23677CFD026EF853B375D7AED73CD54A7EA6577AD37202518963E4FF477248DCD2A4F8061EDA075B8CC100F0E8072A30CDF67185941FF01B6D9AD70ACA8415B366C0B6016CA341F02CEC9AC38D70EC616EAF835C25AE9D89A664A95FCA334726858E60D56998DF5153973431A8978016FAA23E12AA9A41C7951F994CF49487601D425B0E86E603ACC22EF6677632A840B19EF351946568E09CE7BB6C44A27F4AFEAB6450D731B5EDF3D278137ADEAF518BDEEE74DE850C8193323F3CD4F77E3A4171452584341E9F13D2D7A0E7FC12DB249063C3DCC1BB44D1E985F5D1C8C0CB735F0F8DB9D3E1EFA1CB359ACADD6B1827100594C2F29A51FFFFF96623BF6B486CA27E52143AEC292426B57712BB44CA4FA8B53C112D6DF1B224C8A6FC0616574248550EA7BAC1DD4D16C130E44C76C7A6F66D3A17AD91C2B0250DD5173A3FE65799C38982EAC0BCE3CCE9A3EF1E17BFFAE0E03CED6EF105D1D8F96877A4AA37B9B14FFB0B70A787325AA808B3639AA98E847AC271F997A695CFF92A71F3178BD59D068AC8A54474A25236851486D4CB026B5B8F307FD4C03B17A14FE549D969DFBD8F882E9D15E913AA4145BAD3BE361EDF734B5CF74864253527DD8F571FE397F058D3BDF3AA75B6B78679E4F9F663F430A7052D705938904C7BD913CBA19A23253FB037B367C6E4A1BCB62FD9B0A10F3AA930F24209D6A1908624BA8F17726DB552959A059E9D6199483747FBC8167035682A3E0F4F75BBDAB6D550C8602CD903B1F7EF21D77865E73F41B8C5B05765D6EC1ABBF0761FAD42B6727D0385A1DB00FCF8532EED5C50241AB52EFCB8714C33D9D6693B2DD5FC0426DD7E279C809C6E3E7136FC8B3FAD5655E8C67223D31F34991983210F1A7133F5DE6D9AB2A50DE12752D0D7A6E54D5DF878559F09F1E3937731CDA961C4C00F48DDE2D99CA5CEAB88CF630766976566C3E5E6CF29BA10D7B70940815095B18B59376E0C4C1142DE487E591AC89A9DB8B21D3F124F1946B7E92EEADE83172AE2EA2CA2034F188403F735E96F71F906A2E8C3987B779BB8FB3BBD24D014391331EECB14CF3D857B4B99B7AD071581740DFFFF18974918ADFEFCDF89CB641DBAA53DFFF0E60706A1005BE2932599B4DBC48888EECFDE5130DEB11BD5DE85D72D2CDC46BBF045FD96EDCFF6E879F75E19D1BE0EA2924997EBF9EF35E39DF370F6445C8A83B28599D22B1A3866CA4A201495B9C94F7C1B89B760F9418A1729B12536C1329A0CF4D29B0D8ABD1B01F7E53A7A4D0D4E19A6B876F697778520A75CE936395DAF849A62A207E3F63492804ED87E62317412E75F9471B7356E96DA7E04BE509C50CF639CABC11F36793A292E2C060E5F9FAB1B39D38A2D13214624C23E5C315EC0AD55E6DE01DC8F4CBBE9C184D87C925918DB351C1049A5B5419E88506BF163FCAE07A89967787AE1374A1D2FE355BFCE742D2FC02D0CC755EE4E567CBEC696D819A4DA984B0786489B6329D89F9404981A461701C97CA0889FF3A0EEC115446022BCC3E7EED9158B2FF93CCE9567498F3D17910327B994DD8BC8726093B642D831BE3FE82341B0AC493EBB5E592C51115434A503ED761F62A5E7289E855FCAEA5896FAE6799DC3E21B7F79461B39C4B466F8BF5DA19A6E2CA5B885E723CB2CC385D7981EE0B8091392469E5CA3C41B2ACE4C6AB2224FC2F0B4DB9E82B15529B9DC1C0B37649301D1AAE2AD638B2307433B373D4D8508E0900EFCB1E289B3F63FAA2A7FAA0857620B99EFBA02DFD0ED66BD2736A795D3E35CC7138FC69E9BC164E58D347989C56B72DED2216964A7A39DC3507D4A18DBCDDFA3097074CA40DEBA591EAA836EB1B63A724F8362B38765378759077D551A838F11A32A4000DDC16135D4F0C9DF2BF7CACDD3649B6BDE82CD4970528BA2148F4AE88AAF657C840ED6EAEE403554AEA8DAE5AA91E5656B19C009A6C40EB4AC50760A45788805DC755FB8CA07859F8B730D7F0738F28A998F6012B541F1E3C6A1F173E0C1C8BC27E11D9C1C7EF5CC2C764A97A8D4569EC356CB0D34B0E7F9117B36BFD3B115D60BB5545DD6B6E0659D95C39D3B025FFD60C525F598D3727C3EF453FDE39261F013869A07D2B763E84C63E0A62C26EE64781A5234A1295DA5BC26143A9E2DC87D3CEFC32A67D717B3F9C61EF5782EA2532FF12AAC109DDFD6B002DEE96A5DAF6B5859D5CF791D56A2C662D28100'
			context:   '799FBE4E9E7F32DB58FB7F386273FBAD48AF8901D4651CFE36971FB738FAE2502B2D9FC11BF80907CE5CC58683305925487A51B18B1F6C1960'
			hashalg:   'none'
			signature: 'ED67BB643888E817D22569FC311D29D63EE636385B6965838E49258036E35F93E2CD121AEA3AFEE5C851888D79D2B657AE1FE0CD3F07CBB129B9CB66C5F768C27FE3CFBFA3FBAB24C18FBC48A2A50A8AF27505D19453A5BBA033D1D3566778842A007539D26575CC72E513F8CFE0373CBFB67642DD5B4C838561B20FCDEAE3B897BA4B1C24A2142DB9D98A3868E97725C93EB131C1E4EB3ACA8C7B074048DA52B809C08DEE3E3735E6236A96AB298B707521B8DD3DC81F7D3A73D76D03A9B1451C7E9A64780ED7EA9A3AE8CE3106C55A1730A4A18D1409B6EAB875989A75F30AF70A1F9E944832A1F67C96C5B1123EB4780604566CC73B250177A726BE66CA332B37E6479B99B6129CDF8339D49709106258CCE0AF1C914B2CD574E897125D2654B33A3B2CB77CA7CEFEA1E259B8B89A50E97F4B8148AB684F4B37EBDDF0DCFAA195AD1C40DE51C7498F549571EED58FAB1713B9FAC07230BB8978E0C1DE0F9B7A0D6C1B49D98EDD68E72ACAE97B3E7BCD1034B5DCA0771A62DE9C6E40E10C01FD02E3673954CBD37BD57503230D14FEE247413A8A1EDE6DA14C26893AE1A144AA6F597D800C551B875BEE11B06CFFC85A17F3625241B1302A1337CEA646BD1F8C14B68C1518D934D480BF0C1602920B26B56335D72C9DCFA820EE88E1D1AC368A4D93FAEF6502AFC64109AA586A9CBF3E853E54DC80AB4D264B544834E885C4BBCF65E6F3118FBAECA732218D898F933B5320E632D6F286A89EC9E3F3422E66AE29737BF60A319DA5244610EDCE2ABBE802C7D65C728AB110E9458915BAE878FA30484B54D5EEC6D8FD1BED38FCA537E493B0A126541F34947D734664393B4EEF59C8D5A608699E8F6FB7B3E80AB13F6B8348931404E9911F41230BB1BE57388915634B5E602A2DCF89D1A0509609BA204B083522817236BB511976C2D780CC34E368F27808323F9421F52E84BB361AED00133D25DF7F27352E921FC156642EDB65A174EC02BECF345DCB00CA5F113ECB9CC592A545F7EF39E9B3760255D7252EBD588C7B1B6630145375777306B538D4A7411D986914E90156B1D8B9F219487F38D00FCBA5041CD818A421D030578B11F0EDADA9EFB228130693386BC10BF7BCF3A35C417DF710C3FEC93F0E6375DB90ACD65AE33C61E56C37F7B97C543094ABB2B9911A167CC02BABCB7CF9A81689FCF96FD568A7B7903920E57F90D68EA2DA60B83EAADB91A865739B338F470A8A820D04F76EB6BC08CB7270E9F19CAFC1011A4D375ACCA1E0F77EED621E8D5DA269B6CB22CAB3C80B57FDC4FA01EBCCBBB0FE6186A463D2B09F902B5D2352DF79388FACA0A8DA63D1FF42DE5045BC85BFE7E1E3543089D6F6E201C16104ADD7F5B9FBB071FD67220DC60F30B8E8888A0F998DDA951DD739C60D8F8EA013ABA554F35D9EF6AE867CBF6E5AA1C0E2B267289807940DE274B732FFF562A521000FAF892BA9F2767D9E42409CEF6510B51F79C437EFA9DF5BFBED5694AE7D92CFED1BE31C5974F7A2870D651E9173D88EB9FAD73EF1627392985A4A82E58DA05525F817D45ED52905AE1956FE46FCEEC0ACA2432F44F0F381D847CF1F52F9D208E2586462C650AF28091B21A9A9279381841131A32E0A4D36EAD1526317CDD1AB6C74BBB3E8F3C9936895C1F5BBB080D3705B79DAED2E114D5DB00AD565C4CB7358B1F6EF69C540F85659D780B7786BAAC6CABD828598F61DD4AA4D65FCDEE0392215AB51D0843B03E8DE3E93D4C392AA181A5F80118017C41CC394818686A6FE42085FF5AFB2A7970C901CCBEE168D7448050BE4E5A5591EC69F2ECD26DEE87EBE6AA6BC2C7E683DCE82C6D583989D464BF042FB2C7D72109F2DF3CB897927E7AF4540B87F5DECED1F4CBDCB300EE4194B46BEC0E71641231029375FC3DFC26E0F6D10A4198A5EC6105792DB7897C979A12480CBDD6D19FE0AB7E22B067E6E5E4E2F47FFEBD31F8C7AF64D6185F0D27B0FA2D0C8FFBBCD7E954D389A492F358F350E581741CDDDBB1D098CF81ABAA59C2D4D5251AE6E2D150DAEA3DFB87A546C9E6183183BE639CDD9E4E481121A8BF2D432259A3CB145DCADE90A598654CA9089D7505D2F841902947BD4AB96ED93B0A340F1AA05B8CF7E758096D727F68A57E4BE8D2D1C5BD9BF5D30418D27B5F5689A29A8794FDEFFB03E8CCD8D9BB78DDF9DD56F23F4B6EB653B1AED8B48F03BE04F986F576D64B392D81EA60A00B2FB2CD1F22AB7C46093D17F89A51DD574D4EFDAB9BD57EC5BF673319643DFA4412CAE2DAE3DE55EE3828B3346E13E051FA15906A6125A847BFD006251A704EE3B846D5DED4FB81143BD2754F7554BEB6DA03500469960418CBB3C8613DA7C6C3DE833B2D5966C96AACF7788AFE5B281C43103CE31B9CFA9F4A66060B6F65628BB77AEF5025FF981F09044732BCD82D968740F29CBDC2B0490778FE4EA004F000D2CA342B9AA8BC63508F1DC329F406DFEE3FCCB21AAD6ABAEF60ECDF5F62ECACD267EDFA7A1DE4AC7EC284B07D4D0D90EC9E08F9D8128A0353E0A1AFD7750D8760C882AA8B18197D14D59823EB03F435289A768971FAE3832E0569AD27CFF1813C7A331C4EC302F6AAB6C7C61A79B6FCDEA438D896B3530979A7A7AE1624BA6A2D7CABC0A9B1C22C854EA595EF984DEC064E70A1FA043A9A98135E13B71FF834FF537E78B5329C156A6BA630C87F5DBFF63B16F9A8C34BFBD6CBA8A154ACB0738668ED0E387395DF679DB6DF467E79A06AE55932772559C897C697975E07D79168EF31680ED6D4AEE1A6A52654C9C0ACA3894ACEFAEDF8500B15F00C6790024D91F6716E525ADAF46AEA014736EB0FAFCE6258FDD049AC46B2865C9CA696A67390D2EB5E96645B95F70DF25FACF6DAE822F08F0E196C66BD2C56011BE545838541EA5A23696A316B9B6C50AD92A0FE54067508F28C9BD2C46DC6BC50E6E34909E5BF87C7E8E2B303923679193659A5D2C34941CA2B337F2D0DAD741D8564BAABD84A29E7D4F6A260CAB94F9C3F660056B0FEA13BAA14743ADF31AF7346B1765DAB04786B48D22E8D7E1B9C8249AF107808B40F166ABCB3834175F7BA5C9FF35A775858CF364A484232CB4895DBEC2B569C10A3378FCB0F3C331B0B177E1DE21E4BC10D92D5E233C1F70324097E0790B5C1DC5C6041005A11AD832079D259A3CDAF865A4AB1E8903CAA3F4CBF06263E1EE0804EF68BF2E1B8629BCA7B69C32E59571873C73DFA037B5FA3383335C03BCC2EC181A574BBDC3D7DF3AEF475D073D1366CB9EA48DD63450E43299873ED4FCE981B34A466A1D05F7802131A2278762BA12DB9BC9EBD828FB9E156435568CC6DE4119C280C67C698650A459D51F0509180335D77409A19F6ECF0DCE6CCDD57BD12E60717F69E64A896E920A72F062AC5A2D76FCFCE8F14D1E0B0F622818FE7CE48F0ED1190959E9E137BFB7884D42E0FCF34E961A0654E596022140FC7A751E8BD3BB88665867C2471A00A5881D04570BB5DE6D53F1A395A4C27F44CEF05802EF26E34450932C8B911084265EFEE56E12535C9AF3BAEDFF3FB916A2B88DE054B11173C13A2D22F180C3A7F67110874F0F5FBB16AF2218B53391B7058E887819E829CA7AAA2873ADEA08E120C44EFEF66063833067934B33045BBBABB41F058D8B11CB04EEB6412CDFE107C6814E684C3573BBA0853232DF75ACFEFFE1F440BA988EA19E21432490C654BE910E2733116794CBA6005ED331628A7FD3DC9B2819F82C987DC569255ED2E239FAB3F0C2F3BD3960BFE04F5A0C3B3AD374CF5A1A467E678D3B53FCF8AFB240B6F6AA7731E9CB121EE82765DFFC4B3221F207731B6A142487421BB7249DD450D9C313D6E262913DBFCA8969B118F02FB196C78BE8517CC0D4CE1B7DD18F20B2A31545EA22EF338BE226FF963F7F7F712FE460E43A3A97B54F581476F7DF78B9420F0AC730CC4830C278952117B520396BB6136A5CC378F5C71184A8A8C52EDF79C0F43CF0B4359DDD46D744F0308D50C624B4CBF1B38FA0A1528D7E9A38592578CB1DC0F58495C5996A208C9A5719C72FF36C74DFEF5205C32BE0FDF997C1B5BFF174286D6337C196FF9B761357190B65FA8A0BC0CF1F07EDF8067847DC4E83C7CD8FF0EDFA128AED90B49AED766C47CBA146354A168D49EBEC4B414B16B46A9364E08AE068AF9337E04FA0AD9CFF3A54D4F669BF850F44A5D50B72C840B1D32D6045199153A3457729DAC6ABB718ACAF10B4635A88D8B3D58729F735A8819AE97806AC2183C576366E2BBD151C8728E9E6331730B937A0310008445134F7CDF31AA0DF59A57481B8C453EB1DC4A3EFA04FDEBD2C4F80763242AC6C9B37FFE6BAB00137039E10585E7F67F53A91E00D7736838A9076CDC6E895CA971AD0C7EE7E786C45807ED1812E82DC0B0CE20366890C1C1818EF7FDE941806309297EF445AF9B70A48A414EB4D2B5FF796A1F3CD19FBC4773F0982E37EAF1609ACE8E088587F06240BE88402A4C9C2120533A2E81D6FFDAB5E89B6D57C09507BEAD423A2B65959A1B78441FF09D9DBC9C7C6EED4F1C31D775DF47F9ED1F3BF3A29A93FEBB206CB76430164F42CF8DF18624638DB918298094E3EA5C71D2608347D11D300A15A594CB11804F736DF96BD6F261264C36BC85A556AF85FADB579DA5A773758D6A17557875E74FAD20916611590495841173ED9B6CF110D428FD3C89AC2F945D8AFA92D2ADA44189362EC055D88CB50A262FA738998C1DF500DC8A77820E13D19DD2AF14FBB179E84E936907DDA4B8E0C7CD466B11B46399AD388395103910674C70BC4C2CAD3739D35226937E533F1034E03999959F62AC94A37CDD05C81B7D031810D63FD4139CB1A2681DB5E85363C734C37DE1FA7CC4878D41F3929891E35B461A3CFC25D9A8FD0A94EED634A8862819EC75E94C178C5965C92143CD532C96F57660263137C7FFAEDDAC3F08E060999A4B51DFEC29219CC6CF8802B0E25F1B660CF671D9643B03E6FE0783F21BFF28FF03074CFA93523A46108805A32AA32A915FC2EE3267C9C8353764967C47A862C306BD562246E2DE793A7698F9F31197D51540AFB77F928964CC99044CB6174DECD2235B17C0A8F7569DB32CBA37566E87BAEF2DD840A4902C16D1D051C359A2A0DE9EA4D236434D2AFF5048171620A111B286F2D83BA77547E000F6E41CA59B8927C6F3BEED2F82CFB62465A7A87169FABA9C494154F4C3FCC2308E93456F46EF77D5F64E0EBEEEC24946AD06C950D31BE9B6609822E1C406A1E399CCECFE16285A02938F254C3C68AC7C1A7B698D07B82F2C7B13D0DE5E39DF6C79EC1722889F7F6692645D59386207892448344A93475AFCAE57FC2325DCE666F470D8EF445D64DE7049D9EEE489970EAA1804121EC11A2E28EBB82779598B1D6C42B05FC4F08C7D7867C08EFEA150D525210189AAA1728F91E2EAA70247893470E9D7FAB42C520260364D397C7C35E58DFA4758048B6F2585421024E1A75422594ED374734C8FB3A91AC6737B95AD30C1F3FB12626147DEE18EF6251A4B208C8DB4404C984DDDE0827FEFB8EC67E2FB7A752123BF5CA273FE4484E680E04B1C5C700767B21757DC442759B120E11E1FD26967FD5CA987E72519C989493D8041CD4399620EACF117B4DCD3FF31CFAA810EACE65351D10F28A04C7BB64D5DEB22B147670674C5EA03DCE7EDF2877A47C465B822735CAE1251024BCD7D5B801D6255805DD96DADDFC6B4FBA036AEC3A4029401C3FB279A97436F11DF012E877E766F93473A3FBB5A7DD8EF3A512F437AB275A8E939259080D8E2EB8E5283A27E349DDDFDF9689DC25E42D6C4874D031AA23FCB4D378DB9D7AD9F157C656F4B3EBF581AA9B147BE1FB1DA1B6173CDCF24B7A091FD79CAE8024EEDB9000350004BE17FA36BF72B45D6D60756323A3F67A7FD0FAFF9ACA4C0C3AD425753A1D26A4FA6D806233ECBC5D912A9B1470B1619EFEEA814CCCDEB83EAD964031198D38DB748C973D61EF8940B50AA9B510D635683F110CC079D2D984A107023DEEEAD64127C2A7FD7E9498E17CF268D314B7C506F65919C7BF480B98AC94D131E6917550BD924C30C0126B2FCA9683A445C02A0A3F0AA2336A5E6A2C3745E044342D648DCCEC17B554F7536DCC3C2F4612FCBBD700057158997AE9368217ECB2D7276DBCA3702DE8C20857222C3246F8DA11843223D87B214E8DDF03B82264155398582AF7840BADA350209D79CF303A632DF60AC94EC10A2B8C5F119C1DBFDB78C801E9DEB96ACD8952DE5A7F3A94AA543CD618787ABC9587281AB9196996CDF39E28A368EFDEAC1BDC5B45421D6E766E587DFE1F8A7C23DF9B40E31B7093FB0C2842F865D11A0BE3F85A3812F9C48A1659A8E40924887DE93A12FB96CD07340D90581F214922BADA01FFE8B3A4C4C22431D7F90718B2B6AE9C1988C5217B4895F24ABDBBD484584951A868B3071C03872A4FF15287AAA0F787BD049C4955D721DC5132C301FEA3786F91B07089235E01650D3A0B03E74FE7392CD672D9C2A9834DD3A47C0022224C880C48CFE174CBFCCEC20F367081336582E8D500D97EFA594C22D0BF5929D8F0B1A413738F362EE3F4EF80D688871652AFCF226F164151C777761BCB42FCFDCAEF4C3247BCEDEA2D6F012C13F993D69A9C51D33C31C4005C40007F742BB6A7561CFA5D6331A3A9E95C7D245C1FEAB5FE651300C188E0D4B6E84243925E90468B8F3F5D95B3515EBCB04B18D7C2F5AE64FCF8640E14E364AF483B73DB3B545C4B67588B93E0AA986A0F76867785448B620ECE9F7F6A94E08F776178F763551EA8CB020B416029C9CFCC8FF25390138A233A755A75D60FB297031D77B96BB4E72793128FD16D728A0854880FFC7FFE295E7D4D1A4C65BEC52C818CFEA1076CC7B7DC94329DFA372EDF199815C1017E65126B1488FE7C22D489EE3878F62D5C1AD335D5E5701A24D9CA48059368FD0EE66456252A2A3F38D68BEC945912599DDFEC6FADF7A144664203420EC888A0C27CD75BBE07A10619F34F479803EE43F522145E5DC4BE55DC2ABCD6F3FF8A83C98A1A6628F0906426AB48AD3C0A84E3AE45668E6C0E4297077FF74314F86E44B0A3F50CB525B8EF64D8F12DEF5262E43986D7B070C19002863B1BF50BF0911C8C1F73BA27FCD944A476C53E160E07FB7AAF88B1224456B2DAAE0E7B7668BF8AF9257159563ADB475C5A2365CA640992B90C8AFDDBF5D33153F004E4E09228FFFFDD8844103A6B69D4F27FF93EAA0C86037C1EE2125B86762D43C15DCA709D9970054F2FADED048D8B00D9FB537F03EF1D679104317F62848B709913ECD6C666DD727F36D3DCDBF418B81E1BA6C7B9673F18DC66E154B8EA7D20EA3213DCDD1A2B571D5D5D480FEB5D6F17E4903327F0D5EBEE29A86A2ABC5CE624E101C58FA9B4ADA8B91AAC1D6B11861622814E3E32086F7C5C93E243AB395B041204FBAA68CC477BCADF8939F3FAFC02ED810218DB2F31F678BF44329C878A3DEEBC399B422C2F7B6D596CE275FF7F7EDFD3AF4966A9851D8CFF85095485421576E63DDCB9B0F4A7464BD33691035D398F93C89F9D7B75215447663761307F503B801DAEAFDD0B4FD8BED3FD74640A896ADED13FC613C25E213C5623307568CA481C8B13856CD7542121480295A466B933DD5CD56F86DE97E544D74E4F3E9B92E0D496DA46001C9B8DF641F70E12CBE13EB56F353D9C491CF1F81A7A47A12ACA20433C47DD3FC284729C8EA349BE5DADD88B30512CEFF6334AECE3432AECE4F952B9D8523619818F1AE21FA982C468E718208EE6C7348E591049C89547DC77C4A2207EFB0531F561F0669752909AE686E2E34422BCC86D93146A5651DAEB19C437C7A9DC03E77279F40B906BC3E1DD526AA7AD6D549A007A3403A266A69A7251DFFAE5C39EDA7D242A329FAB6A00FE1548B02513F0B846F9D6E1919BC6A2E26E33D33CE9D7442A005928C48044DA40D1154F52A0E8E496DC657B0E18E22A3847375AE368D2BFE69B1A63D1D35C3814CDAE339E8C75BBD18E822EDFD364C1A4417D73BD40D3A2C656FD96235CB191C7081CD1855A6DE69CE97B432D0B1B2A94A2ABDE203D8BD202C4667B94AA7CECD3DC63916815AA9B3A501A65B4952F3DBB114AC926CFB34CB508A7B72E00919B91DC5E93A6C5B88B677E19C434BF44CB5583E784AE6D5BF62D0D8CA03A41927AFAD400EDC311BD9D993241B72280CDB90D711475ED360576699090E38F30280CA3132561A4D7264C3370C47CE3BD516502CBBEDED93F4A4FD3C8C67A5D56B251522A2744FCE84A46A4EF3A3C82E445DDFB335FB6E0A181E6EC0D5D78B7DAF75BF682CE46BAB1FC8562F1E1882F3598038851FC6859F66093E1FD115A9632D3B063E1101F9F46676DDD15541A9F3F4E7A20B39FEA99797CA2B293977990DC5A60CF46A9F6AF4E24522FE75A8F4B2227BFCBA79413448EDB9B1B2EEED308AF06AD8F28C6930AA8FFB834A19F3A54A749BD73C405C95F7009694212DEA83609277930977CECDFDE149D227501D52A83806828056AF1C90B5EFCC6EA6E3E2F4B7FA90FA2D6E65CCB0FF8765BB5D473CAADB00FBFDDB71E08ACF8A900B383238BC5CC4C836C319569A9BCFEF3D68A98DA16DABBFB2592DBD1B85FBE2F0FC4EE17BF166A6DB7A4841A46F204DB82A568E98E2A5EC207AF7FA3C95DFF8A8FD608E70ACAC0FD772620B00167D84FF8C267D1ACE08A88302A6B9FC643FFD097E77368DBEE1A492B368B8346BAD9DA43C0337B41ED966394A955B441344AEA0A727AB97CAB9780C816BA85808B93A945A8F53B4F15041CA62041710F0215BBDF1EE73E0DFEEDD4C8EA91EBE39A1F60F7A66460763EAA3FA33C3FBA3202A282A35D43568F76B814883DF33E4745C07BAA1A7485BB67F6E43866AB403946C8753A15E2FB0D3716C78F697EB282A4E28A65BFF95A009483797FC0767DD4BF44D8BDE48CFA9336533CD6B6EBD4B8ED2329B6402FB22FC7FDAF7AE7C11140F120B123227004579E2E7D54D979BED0052CC4534DAD05007589D00C4CD885D73287276759295F79333EC420293D6C90B17ECAC1E0C2F2F8A8E05D23D9E11B93B31C90B0150DD2AAB8F2FFCB1152490F11E0CEED0F76A6773966CC77D99265FD602D76FE462E0EF7C78E7897E8839C875D8EC867AE66A166E831A2618FCB8816D83F804F8ECFDA5D08EA017D2A0D5B571F914A2831FC2235D932759DA753A6694201256D2F6EA8A330B681C737C29B8A7A0244B7760CC435F2EB250E8000940160AE91CEC820A8022BFB41A425B2CF6DCDA3728D153A22234ADBC4ADF46FAD7CD7B4A80700DAE87A122FC9D18A54052BACD1A370A699F161004A73EF8D076DCAF70E63174106C7E944FB57A7F82534F1EB37B556041088B3DD08BB5E1B9660014FD045A3F027D0B508A53FE45BA3688078B97E95A0FB8EE6DD2C1E00F06F2C25B5FA9054C09C9DDBFC1168E62EEB7E76FC2FE262B105938B964312C08F1158653C35A08A9F367E486E1504EABEDFA9E6359801A070DD6B67A80AF7B129E1EF1F438151E3965F706199BBB7717264B6178BB2EE62FC66ECC532E0A4247769D78AD7ED98E2155FFE36E095BD87379CD825951077AD3E3B947B71240D21C885C5CC0F2FD9EE9F050318A991B5F45ADF27684F6765D615308BD343234D0CB55BED0E400171D03A7B2FEDF4653BAED0E350925A3241DAA1033B90A4A2C074E405C0CC1DC6E9C4A5F701462931971F52BE881277AE3168072F1FCC92E45D0F360ECCC2AFA8B0A495F19A0C506BA2BDD62C3E4935B63ACDA17E8ED66547D71EAD4F0CD610FC0E300D97AC67C1870CD0CEA5782DA3A249F4C2AF7C88ED25918D9C5B6ADC698F13072F6302DAD0A2266236CF8D4C04827C10A13E58A48DE9E3E60FBEBF2790C5FCD43AD9CD9360D9B8379B9BC28CAF2A58147BCF72BAA94562D77AFC2E2591190862BE016D239E7C49C46F9D386CAF2AFA67732AF731A4A370B216F3B437F1C12D04A6740A915726A9318B17AE871EBEA667BCB999411735DFEC7D2069AAC4E02B5751E77BC8FF10FF61C1B74C88F5B9D4137F9D49BDB45236F5F31DB5C33EE771D9B5E95D76334F69F7FDED2BC008DDF7AB3971AC9CBA3F6A09D4EE84680D5760F42E6F9C5972E63B01FBD518043CB06F0AF858B8507C1C34363FA3570FCB1C283B5D92B38218C74763CCED43C5237503472861DBA0173DC9683894AC372A25A0C73B4491EBC2ED3D7DDA1A667B4C4B2CA4BC433A2F4ACD2463B354B52EC642BDB887F037067DD2D1976000E30FCB958E198FB547F380CB6233E3EE899FE82EB4427850D48CF917101199EE64ED7727F8509585DE58D7CF577000CF02378277CA01FBAE65C4263E4D51F18A6D4578FD47CF2589C2441092A4BA3B9D36570599C213B6F1A0EBB85A1F8CB682766D8BF8A2E16D23E7527E5985A726E35EEB363037A9E7AAEF33D1D579D6A7DA434B2E7D5374EC06A14546500E93845A74DBB95988897D7AEE99143EABFFF5C1087419E9CAF1335B64301917EEE645D944ADA2B511B66C15B973F27A385AAA4023CAFD2C2265CE2DDECF09C0669314EF7BB61C3226D6A1764578F7CFC771531D8B2A5C289205805B99E0AD22F3C1A3E6D2BE2A8D9A397294288B3960D16A3D31C5CD22101FF910757C3CD6DE94FD1A19B17E6294E9DA00CBCDA7FAD7C6FC7240D30B0784F5F369D2FDA1F9973B29273DC317CE2200763A3C8BE0C016A598C18641857C45A092D9118DE4ADA25286C038DD7B48EDDB30FF4683F96EB2A95D1B3193194AF429D813D6DEB6FACD47507058F58EA81A520D5FE4130786EC1C7ECE36D499E07AA1C930F8685DB937DDBF80BFE9FBDBEAD9804EF7C8D9F3506DD79461D2359FB686C5D54CB049C4A036788B8C3212E7091BDC0B24885CB569A9003636946AB239D9D1C9404F4AB2887DBB7388BAA16BEF8759B0D0D528590345DF95668A9D50C9A6BC7F4F2CC018C818F1EAF629CDD9B7DB65B0059FE71B8F5BF41F7A13D19C5E61002B4CE56AD85214FC1F3E8E7355F4551CE8BB47B104F9060B1AB81A57566EC443CC5236AB6521BFAB1D2F8A502C6044BFDF4904CBC0473169B2B25B2861AC267BDF3EA02520224011D9E1EC23F1E62744B16C50668CAC0CAB38E88635215F71C89C556993DE0C2796B7339D09A78A1670B8738445863628B6F1F2954CCC56EB50535CE6CB8C57451C125433A959117DEAD1B3980CF412B4B3BBCCCFC8FF771771EC18FC47293A6E80AEF96333BF0D0292FBD3F46FB6D4624AD6B617BB026E1D8F3B2F8FCF92D3351B31A2EA5E9F59D96B13C15803D7B857996CC5FB6B17FD00E75F888DCC3FA18A5C6513589B7317A09AE0458699FAB498D4EABBB34B720853CF609031FC48C4FA78D72DB88FC669B46494DCB95B2EF0161CE3E9AAAD1C22D710BCFDD491CC04DC5ED68B6C51C9182009866F4C95922F771F13B800C4E8FCA95E8FB3A0E7D45016F33584F77E4E9D90960A096D1FC90C9F6B398D5AA8035CAA5E56C4263AE39936A84BF08D59AADA27802E1E877FC522D4E7149429EB6F73E57EA5535060CCDD376EF530124DEF977285C0BCDC87F1DFB807216872CB3670E326CA5170C461BCDDBF780851A06A5BBFB67C34E1138639AD32D9CBDC4FA7BBC981462141F39EC6C0903B681A0CCDB98983A0894B1A0923D8A8B172CA3E8EC3C4EB7D2CBECE7CA93CF607E5FA4300684A6D24086138B3D6394C5A05318FE088F51F97406D7F6A8147E44A7AA0AC8EE6B223BE4213AA17363D55DA647C1D67D54A52B7D4E204ED36BA9CD722E8B6183B56030311522BA076D72D5C0133B0F56EF803DAD8F58198EB6721DC8C0F7EBFEE212BC024A200F756992E8BD2E9B1B1243F3E75DA2880EBEF69E73FB3982D83128D4298153437E179EF166C0EE600B1D00971523BC4D6DDE8D5DEEDAC47B94DD528001FAF02B9F43DF5E41CD4A925DC83BD9362F0D94A64DA672525A82ECF2714A917E7BED23F19572CA846D8ACE94E9442C72AE3DF9E14FCA531AF64F5D31064B99FA6BF0704AA0258F86624A32B7BC93C8D0EEAA41483B2F2DABF2B8E492D4CD07D57FA39DD90788383B6C063ADA1834A8CDAD0A4CEA2FEC33CA4CF457ACC94E75DFA2A0AB71A9552B1712A2137FD2B9D3D444678433FC89BAF6727CA8F2EB0617B73CB2379DE5C2CA243990627C224FD79A63B7190FDC764130A8A32D5173AD6253F1A665C7BE1CE6620452635736F4B2BDC71CEBEE747AE3382EA92721AAEAB8D947DE8CB26D9B45FC8AC41714754C32C7C0CC5B769EE3FCAC6E590F2D1E16385DFCD00B9D2FB4F3FF2AF3B2062E7FBC523F149E19DD25F8DDE36F232A00D5E90E32D8ED5C636F7D0A774D7C1578E25084FC93A505DCF90030FA98A35619D96408F41A5BEED296063FDA91D6B681784FF7A75CD0EB0E217E2202C9CE2E4E4602B337A79018299737ECB5FB9A7C196F36C16BB8485A81094DBA7CC054501113FA94C8C80EEAF3AC94AC4A9303B5566A7FE837CF4EB8EA2335061A1D283FC426B8B948D4EAED7B6065D87C7B06ACAA84F4BDBF0491E0E3D96518E04AD7B66D5B774DC9D92908391200F0991BD7785383D2DB50D294D17A655863AE13734C75184EE4F0E9AA89561C673B0638687A5A1A98EFF38FA950AAAAA5075B312B6F5EBCDAAD3F21E2D64377653775767E4B5CC56911CEF11E7E93A3943A81CE34CD095714918F637AC2FCFA4A44B73C1CA05F50EF50CDAB1FCBC30E5C21E379F4A38CB34CF86FBEAE60E369D82679236039922DF47E36F882C9F8222269144AD0D50463653FB5114CE0E7A6CB5657C8E8AE8EFF1ADB3FC0C8359A86E211970725C6B537DB3990C9B9193FB03FC0F23BF07B9B45C3E44BFBDB7CCB085FF2C9771A3E3E75EA8946E7E0946B675F4AE5784D041F88FDDE2DAC88F0DEC571C8BB024FFD972311644AE03A7A4B5ABDAFDE4A6BB2286B66BE3B63A1E7A8369678A66257CF9413D904DF5A72F2E560D84C27F83592B3538888A85645B1E03246CB14BC6BFD423F1AC31ED2FBA23258FEC006147AF78D993B5D6624056892399FEB92D27A219C4950A05F3C38320EC861A19BE17707094A5E5549DB5EE5D42AFBCEC10F91D589C9B3E5D324A8CEAB12A0DE695D770C88DE10B79AEF23DD3FDE34C541BD5D89A8D2170C326A87AB6B33508297BE2B0A246C32BCD289DE1725F6E9D6855559224FD76773888F7708158C9AA8F8449333FD4997053DA9D69BEFFA540D76FC6B4218CDE30BA5C7912CD767B68426B574F2638037191853E7EC07295FC36396A17648A137CB289A415B6C16AEAF07CBAE18465BD10AD4758D908026E3DD0A560384883F790406A9395A062AB8B8D284B570569B59B661A86987B8F701D93D41D613BC0F2A86E6928D3616FB94F67163A1F1E3CE44C333B870B8D0B5260A20DCA37F4EBDC53B14C21B5C104AD148793C9C8F6EF6B88C0E16F7E90B01E2405E41D8B852FAEF3AC60642B4989B523809F30CB2A179098B0B93E8147F00EBF4A57E87C4CADE2656FBE000FD1AE3BF257F977D44EA0999BF6B4E8285C22DA016CF1FC8BC71968B311541A2006298EAC531467BED1BCFC1BF4358331D56F9B1DCC311E12B63F07F43A0931C41A1C1D49477B3C314AC9D79BEF8B12C026404E204D3158B045D265FB353B5474D7E4D15E5C11D39A896DCCC7EBB1F9CB38A24DDE92663E427B5EDEB83D58DF417CB30E9843CA8582016F4015D478718C453F7E4D71EC951539FEE1294EB77327810AF83E421490F20F4201E276B39996C8A0A3727B574AFCDBF46BABAE4C57E7BFED63DDD9D08184A99EA30E88CBE27B6287D91F55D71C5F5D68A7749832180E82BE6801D57379F181896C959672D6D76373A79DA883BD20329799E7AD54545D3962E8D12872CB9B195C4CBDA29BBED6657284D9318512EBA4EE87D381749A4427BA6FCB26381496C46831DEA17D53C625A911CDD48194D743AA8C1CDE51FA8CEA787FF3B5479EFC748B62DC5A15E7F1B1138BC265A7310CF970E4D4701D0DF9E202C6AD580D8CA2C121A30628F2735305FEE6307560E536F09B6F278543B24D848631938299C29A00EE82226640CF6AF81B0D7CB314917DF8A38C4D1B263E8880965F49B1ABF5AF9C0E602969A9F0C2376BC775F06E50E287554892DAB570117E83039904FD3BA05A34CBA49AB14BA29D3026EEA130670942338DBB5209237BD28A5355CAE08FE2760BCAD61E45E0E1235D11FFFF54C7C7E0DBCA6B6D0688E3E564A9AB2AF20CD8C1FEA028C464A8A4DC010879A36E741B5FEA0E157F85C187ED2DF3A42F1642EA328DB861908E9749BE01D15281A4E5A93A81A1F3ACFBD5E6B23C3B4C7D37CBB572246081AFD19C581E63D190DF9451116C127F1B035F0B54DFBA8BF2AF01B43B43AE238CCE1D79348FDDEA5A5D2E125540A24C956828136A6270A6D97D79EA726232257FAEAE33D74693BB977E328D52BBE289940849A9663D3074DFD1C809CE3E243FFABF836B5BD0ECB49B7661199E65C6DF6175D7A0D879E5F554681299F80250E8640C5B52CA607D8C2308D20FC76DA3DD116BD14539E414ED7924DAB85C4E619AF040B026B64A3502287374B498AA2127EE9E15A7ECA9E083760EDDB512479E9703C062F18DB7989CFFFCDC19CA2C95C8F9244E5F379DC6221F3AF32C2FB4D712E6A3FC9B8E96143F7FC55580458B3795C400AA38DBCE57D108C50F6DBB9A10CB4F6DC99C877860B435F0F0FB87EC95AC35CB8DC51524833E2652D7F86EB268B56F12BA4C450DFBF6066A322CC8861AAA1108E2B4308DF35A3031FD16CF65D256EB06A3377B9A2026329E1ADF444D51518395BE240B5D2B4880A030D01390212BA40EC9C1C4CBE5E048F9F59BAE0C9DFA0B27BAA544DDB20994AEB87B595B221C56A822C5A1DBF7FC27DB21E04B531CD7B21E6CBBB10442DC52FB8E95719CF999315301C0F052D7906A0A695D529BCA448411DB6F22305EEAFCC3D79C850D1D7E50423E1932672C355F3D5A13905193735F617F7A27C362B18C1E35E33E5D55E4448CA336E09E77ADAEED2ACB706B5BD284451CED67737B69364616E556E251CCC825937751FB5FC30042994F6FCBD9EA4B5C71123E4EF3AE261E1508EF8CC1CAD9703C2E6460FAABE90534ACCD817687A8EC879DB573D3C3E64403D4194A4A87959CE45D2EBC1A51168A12CFD7E729CA07C5290805443DDCFE18441D5EC05590549B883E9C6811F9A84ABFDACF0C1A1A2991239FDEC47B20840E3D0417494F26F2871FC780E6FBBD4C8680058991903E9A1B46FEB617ECFD62D8985F0B87477110FE978512A8C65CFA0B051118BCBAD50EB97353775C0544E3B729385421F2CB072CB2A75F33033C9EB00EA123020C8A8F5F5669BF51379F4E1D1589A804DCE0894D45279FE3A8E99BADF706AFB8C40C1CD75DAA59037A6A895376F11EA89CB74BA5D35E22F90EE712061AD425AB28F06F9923C15D133FEB3FEA70DA75A65CB9BA6C867AB3DE98F74042D48D823923233BFB98D2CE2D000B28C91DB4075CFC461614523C42C8FE457054A82FA5608908B3CA13A38D7E9D6372F66BA791A76FB73EB2C7782D653B05E15D4A28D651B4D8EC9F84350AE54848DAD7BDD51AA79F84FBE9FC6376582A68AEC43679C7D81A6229B346E7FB488D4969C8F075B15885F0E49D707132AB2A4A60CD4BFBF5B0DF2F5916D2EAD42CA16BFA1BD57973B512B0B573190058023F1C4F33EC47CD4540D088795B2CB64AC12770C79D62A63FD4D6283EDD698E5F961CB8CACB5537FDE03C439CA167D4B7D9797E4B46A3E2EB92B471805BCC23B8E51E26B2917C19DF2D87B1481592799BF2046DF4052D12C4638CE1257D00CF3245DAF0FFC61A02414643A415D2DEC835E03EE5B7E1158414CA51137FB02F07FF0D8EE8AC5DF150F2630EFBF871B1B86E04FCD54DC6599330D03DE2308804C332CD029AC59EC33409BA626E8758CDF6B994033C72340D12F2D3A015439731040BC11766741DEA479BA4F69B150C700AD0575B033022845BE1175729C8E5C571C15BEFB2D170A3D8234EE3706AB23AFA5124331E9926CC2A4433F403FDAD1AFCB4B85AEECE9F991C2E0F51F72267D69BCBEAC262A5C4D2CE49BF4B4BACA0AC155E27FB8E1BBCB7F801A776247E0C3258A8F8BE7C4C82C53C1D517B69D54BACA5F33CD0E11C145DA7FE371BF38753505DD027B99CF55DD13D98899E928A9A7D055AB4F31FEF6A8742166DD89870CA856201D9CDE8B6D90C44BB1269E395BCC98A21CC69C95FFB31A6BCDCE34C3CA440035B1B428DFBFC6679A222E84F73C54E200A6D12BC338FC3D69691236912E28E65137B69A91CD1F3B1765A6B8EB76FCB17F9D5C89EC9CE02295FBBE3E162B24DF53AE115E4BCC264B22DFCB712623AE1B18B9FC8DA4C591D2DDDF54025C4BCE94AD74ED6F6D68AD7F3D94CFEA1F7B8D5FE8D2CDDBC6496E47EB45F17AA39075136566C91DF435D488644C5CA486CF092C51E4B0E7A8DBF4B54661DA63C6E34777B655CC8FE950168280005ED2FCEBF2C59B54C91AEB3BD522039D1E21704E52376494F845EF1FC405778F7875C4E185B71778C2BCC0994B2D53DEC85D902A38329CD22C0BDFD5AECCD8F044602669675EF4D39BE7DB33AA74C1427448A8A3887ADE6A3C86DB46A4D76026B57595EBEE6BF03BE103972DD92CB36500B2E112F909328531CE7F3623F0D646A28F15CCA9957E30403B303FC302CCA28EDA52F6B96C03AFE6FB9203ED5431FCFF4090405C283625DDB14AB585984CC303265CFCB9FFB045468BDCECE8013ED4DC9E60BBA1734723FC103233651E5D21BDE1247F541C3D936CE14BF2FF50D64CA24CEF3BD3BABD32D1BB18284456B9E33442413893F027B238DEFFDDBA2C20F1F0A0410027BFC196FD7CBC5FBBDAE7DCEDCEBF1EE6FF8C31556824CB16A776C04991FBF039B90DF95BDAE1020E0C7A28612901F66F12B2DE2F8003395A585D88B97E3FA8BF455539A2D6AB9E2767A14E448C33F2079EDA61D21C6DC41B3509E548A714A5223DC6395FE639A4D042F972E281E3FF5D132B875C9BB787BB8F7B5D03B09FEC5AB6CF662ADF95ECA5E3FA631CA2F46843CE77CD036B548C2DAFDA12BBEF917C2E15D38C2AB8FCD6ADFAEB2ABC5479BFF7A59C92E89BE8022DB85042271B2DBE8C91E8AEA2DB678D2A93726A1589643BF33C6F550481765D251B276C8D4E57DB6664BBB9F9B52A082A01F4FE84740148E7E8336BCB24024D35999DF088BD018D54822B1CEA36EC673771C036BBCC3E5D23859B51648C4A53AD132F60F8FEAA72FB6816E2D38A0E35F20F5BF75D8358C45B07785771E694DEC1F04EEA78FA78B6A21E2F93610B3DB4DCF76829E17F5B6C405501783209F3709F5A6F83D5EB88B1B7CC18F883C727C5322FC8C161EB71646C2C0C205CFAAB3BCDD120BB9D335E81CC755D77344F50DD35313C05674B43681BE083B506304DA1BAED4225A00E4FBB35E864C7F649058E67BCD2C82B79250BD22A1407D036AA1B744F0D176F0538D8BBB29D138D7C0E37C92EF9F5201CEF6D8D3359EF8B1819C2933E09AF234DC50E5E8FB3BD01494BE049ED61517514E9895EB1A49FE267C992184C7FF91A339D92B4AD59F4450324229BF1EF185998EEBB4A010C1A9E876AF06F7F05D893770290EA5C8BFF14DCF990CD2EDE9FD99FA01BC87DC9131D1DF29D819BD49D58AE9B4ABBECDD5FAC117AA527EF30C2C380C93A71C938359C6480D7F038113C880DAFDCE54CFEC6BBDEA2D3656D4FC44FF876BA1E907F6727C6170B4F928F1D5CF1C56CA558DE79E60EC89AAA442959413E96B9AD9249CDA6CD4CD1E419E9C319EDD5199C6E1DCBED607C489141284C0AA1BA590F675F667F231C0D9569F672C14FDCCC1E3E79689E207D35ED19B553A1B25EA187D6C4AC115318C893F9381662F29C4C56973EA4DC610F8DD826E8FBDF3B1BC5C628797E60B3A39AA901807682B25AA316D1B4455F742B643A5F68C6A42692549EEECD271DA42893123B4AF6EEE33A44D3E673FD9825280F8A64D9113366CC095C00D1774710257FBF30039271E088C821837C77CBF41DDCCB2CC34B4B35CD42BEFE9B329E47FB188E711DE6AC6DD408C0140316E738B9F0E337BAB2935BB3AF8653B5777A706BC967A52F3F7AD455D6342DCB4F1DC38F32BB2746AEA42BA7AE1ABC1F4405BB58BBDACE8D65E02102916E507D35D49A4B73559F5389A5E49DA02C46C1C81FEF279D0191F0B58693914ABCAFC80BDD74EDB03039ECF9BC80F1E19FDFDB5638419BB849D782633CF5C037360B99F7F13B0AAA33E65E2B69C44B06BBADB5A314DCFAC93A440A6C16B030F5717C2C621C10FECA299BB3920906AE164DC2A1B6AC736DE75D1CFF797540E66950551A51AA72F7C2CFADFB0AAF7640E364C877D40F3935937B76B864518CE0B2224F6053483B87AF55B3F4262D775969AA3AFCD681FA1ADBFE062FC7BEA723180EBCC2D4D1FAA314F2059883DD85683B2C9ED6BD1AEDB8062C0B325471CC061CFBBBA265EF4F94280ABFA255A51BCE090F723D4AA6406E84F46F6DC557063D481B7C694949E6AEB9EFD81BBBECC374C4F0AAC40215064F01762B33435D7B9240228AE13E22BDEE0D9B694DEB66F83C4F2FC6025224C6B38B64A1ED3581C4C4DB5349FE82BAEDD047EF7B46739A41E672DF5FCF46BBC39FBF8E92D2C37C3DF6BA339D4429BE02652B3DAA2FB0B07DB4C39FC837655E3194521F3B57B2327B1E32E4B37430D90079098E5EA60067B6763D79488EDAB4C21726D9AE719E1377E90325933958AF45FE7063DA9129FC131890662DFF1FF591D8139239A5A3A95F730762FDCE81212ABF19F87F98B0EB4684C2FFA640CC4473AB0B6AF862E017B26D35B640C1B46EF58148E11883FEBDAE91E8CA3EF703C2D7CFC78FA106D05295A57561A7AC13F5A7708178E80CCCFB5629363D00D355456F6195AA941A5559078B947C70A30CD83FE2B2E7143564B20E986EE76DC2841AADFA4077C51E0B7C10CB61311F4D070C9E75E642B850075D9F84ED839DF3FF2AA3CA6366FC344DE8772F02277E47909585F7DAF95E72D5FDC729162F5882ADCA783EB30383701436901D6028AE7ECF8375CD9D3DD24BF576365062CBE06DE2B9084D719665C31689FBB3451A5C168BA8688C5F20956A240C6E7E068DF3A2E35DDD8F14F8FD36AD285C86342A2996124A57ACAF92AC89D5F9A3CD5592D491D1F1E4CCABCC2886C1C8209FF356929FBE70968B79CE11972034BBF652BD8D0B399CDD78A0DE00CEFE94F6146557A7E846CBE9260E511F81A489E97F3A4D5532AB222FBB6F32512B5AB5FE19D789240C7A69918283BA6C33D36F5C11AEB6842CCFA0C9511A91C5E80829C821EDDF548627D194C34915FC8C093C5012A3F048FCD9F74550B0D82659C543882F314AD5CB62DA82F3AFFAFFEB081D9878ABBFD18A448E1C22EB7779C32C4F6372BC58A70EF6DACC969BE34CB56B567DF92E4BB198042F6626574B00257C92A7CCA94F33BF7F4621AE25877BD3329079CE401238F2660BC3C5B23D24306E549BA2AC0AB2BA7D03AE500740E7FF6BD8A77D6689ED2E3E906F1D80C5A601CEF55298C354BDC590EAF1D8123E54F35C16B2941C0ACCC067A1405D76656845A6B421CBDBDE839AC6639E9074B39A06AF82436E6FE9BC30E3067A5C1B4B8813DD71522FCC123D7B40518C09F3A94B61AFA9F098939F0942D23EE388A2BA36B7573680899F5CC17659E4446CECE85E47527F86DC3499752754BDE64D174912C7FB4AC5AD26C466623DCA7729AC0295A0E344DC0D10E2FBDD3C926BDBF9F3413F4B688A5A0A94765F634042CFBBD19FF337809F69B4DB9567A1BE9716B7FC76B0CBF2F8002863EF1B3D0E511FB45B075A573C550AF5D30A571529D75A690ABB807814E04E9CE1645B394647F16FC96576255A58157DE1AF69D35F5EE26511A49FB5DE845183A175BD7599CDE390D656805B9C07FFF669667F1B0F6EE15505312E5ECC1DDEF1B2745958DCEBB28E0D1146F031F1519C9DDD6FFACD0E0CE32A0CD07CAA1FCA6F615A7FF3DF763FE4453DA1BDB9AAE659E5053651B421C7A533E4C423E78313EB6E82B83E92BE5ED043EEC3B71404BD521B6B4DFEEA8E709A6C4279958FE5D64793F38EC3B39114393CBEC192D91142AF431439CFACA4BBE2B3FFB8674A97FD5F6A3647BFDC7157B872F2D6F054117A37BF86F2CFF1B1B2ECA12859C8E671122688D4B81853746B54EFFA40EFE49D294FCC0C13462CB9E648C506B86ED925DF2066F03690FA123E34620F271EC372B2440F3E179065A277F1F1A15CC836B8C00F2E938D6A90CDD71C9D7010BAEC02996A2E1B5E244284BE30669930BE3536B98EE1947C922D9629B6235DB74FBEA9B83DCB463829179BFD4EDD583C1C532B09BB3030769802D943559D2B79E67BC53428F10ACC7D54027A15F325A4083DAD4797D3C0CA0C9EE7DDD1B3BA312CB315A39E07DE4603AF27707674E326DCA632403825F871A5D54FC969DAFF50117601A1CD3F820C99DA8F61E012A40052BA8454092F7CB50FC7E553D5FC86095BAA254042451658417F797A81D7C68735ED940215CF22CFD3C0A3864D339C031E201651695AE38BF40C4F486F5E8E9584DAFBACE83055EB6C2B4B4818C05C4A41CC28B8E41DC4A8E98BFFB568B3485C839A111AB7135A7012D1E98512FB38E2758A636DAC61370EEC09DAE0CCE0C1AB398C7BA34D8A833B83C76978A2C0A7C58BAA95D456056DA55BF11AC21AE4C42E14D871C61A6EBDC3247AF0B686E48767D323C2F8B6D96F433335DA5A9E1316D7281C2C08ED31069EB1F881E6A91EF29E1DDF1A5281818ACB5F70476CFBE9B058B8E53B1D7C04F05683B6B47CF5EA2EBCC2FF7F9A75AABA8E5F3A892C9BA5B1942212C3AE185CCCE3BB562748AE97F4EAC45F419069DD62049635F4B049E550973F2414D1F79C4F2B366DBC36753FD0B3B24D251F14501928908774472B10B22D7863C69D59278E056ACE0A3D25B64A31379A8FCB105FE3275073A34E8A105D53FBFB663D33D320C83D003FAEA3312D0E0DC807B58D8DAE3D5C9071A7D2FBF6B9B5762241421562CC28FA2C34FAAFB8D89AB2F4D25712771D2DC54E2197E68BAEF03AF403874C9C606615F155E001D8AC47823FD9B56B2127DFAD45486757A0D9193291E5C51A9FBFD7A9F2980AA80157DC124C95DCFE023C5C7956893843FAB7AAB098D881669D1A352585C84FC06F06A19657179E0C4EE514E79EDAA222364A77AD626227B41F36D541990E83E051EA4F44CF2BD5B7E4A9621F7D25577ED210304B49D8B3A989A914BE6C9BB47E9DE7E31A8CB3B6D814643F61EAD39B12DE82F3C6F28E50C44B9D0FF326BBDC4FB59DBA6B2BC57D41C83AD5B2BCDBC9D2EA2489BA84A25149CFDD24B5DAC35206DC4279E179C2284F5981112BF1064E29336BB8898469BFD7BC40D301D96F9CD73EA1DE2545ABF37535EAE1A5AF672A6EFF927C134318E3BDBBF9DDDB60E02314836238FEEBC049AFE0B7654E2F6F95F1A5C18FE76AEA66638E42D4850AF268760BB5267018D7A3A9492A0BFDB06F4730ADF8087282E20B8B08C1C1F885759ABF0235339F258DB0E27A74A64EBB74A0D0BC531A1D47702139C4BD2B537F645E346C4A15DF008EE00D246F4629BED5D5EC7BB3B8321F114E99FFA0254D7E740CD82E7B000C9E8F0D04486E60B5F26FCC44ECDD164C4041A9E83EA9A1E09EBAE5AFE5B3F6361EF0E7EA9DA1F10B193C5317F7D7D35EB5DD1A58E51FD26948AE28967EF067D54A68E846BAAAA8F8B8B747B642BD48EDD78709827186C5C4F357B9E93DFC89BAEFAB2335A84F6FB3CF2507818193F2ABAF94904CC7EE37BCF163FF5B4A93A58BE7442F3319951A16E585E1CFECBC5766BE8239ECD6D56C765CC75AE14F1A231A6BDB1C48C79FCBD77A1412A6BA6BA2CD52453196503BE8AC6E4CF1E44D621C61F1DE3A686989B601676A5AFE17E0C6C25ECE51D26848974BB70B882D257525DA1B4CB945D33A55508B9087E224E403091FB7272DDEE7DFFBB81262E2DB00028E935FAEE5B25CC1A58BB24523B64516E386232C667EF19B71319432E217028A43BBF8493FB080C2DE55E1D8DABC20F33059FD367145BE50DB9083D3A4F5D09D63E6BE1541FFC96DA8DD370B0DAF0B3F81656E2D27422206DFC1DA08FB38B520403998E3029CB92599EA61A0FDCF7EDE240266797F58BE7AF1AB3CB80C094D1BEC2352BC05A2210216854FE1233F7BBE6C075CA375703A42AA6060348B9D59236DB05F2EAD0473D340E7007BFF0AA68B4EE26CE595456A504201AD264FE6BF755E43BAE2E0B48914B621FEE45BED2366AA2F61315666576A4BB09751DE0BF15B01B6CCC53F16853E798804DE8402F5547045BD4CD3C9B4414C481BFCCFD2190BE2B69D2EEA66DF6884B95883EDA84CD1CF7ABC97875CFCB9C08802A2AB1E389D854DB16D570DFDEA5AAFDFC015D79CFC9B8D049E562A4E4B8168C573CC820328D36990C0973933966290C375A5598F3602B32C67DA07300618292007A4D9FE224E99B3C84B50CF1E56CE1554C5677E0D48FB3705CAC6D2A8945CD127EBBB595AA2F7ACDF3FDD5AFB20BFD8BF7CA0249295098790CE97C0AC6CB6296E6BE0A3B2847E0C15B3B14CBA6F2EEFA015838888480EDBB23156E1DE8669D3560C84C72FC30C3646661C25968EA4E77E538806F5395B40EC0699C43CA2EC00BABB71F1A22013E29BA7315D6B167B2E0057BF22ADBFC8F32955690E8ADA55AC6FE275A57236F4039042FD2411B3F464FF4F3D7063A3836E7D6CDC1680E08EEB393D58E82BBBD05E30898A5E99C9079A59495EBCB26C6527021AA03293A0CC9DC6A41B1AE2AE854488AB8BC55A911C73530B20848910E5ECFBFD90BF73022AAEFF0B1E70D0EB158703F4081643153BBD2B6748EFDE75673F2B0E4430114EBB8E1B2C40683C1B1CC4E28E026B26FB1A766B3F041778F5C69A4388288A6CC088391C7CCB904C5AC3D0DC3DE39989108F933D0C60ADA2906A62CBE7709EC8254E6A033ED6F749BB5DBB13C31AAFC2D9D8671C68FD5D685F17E325F7D5C551BC58705C93B001C695D73BBCE26AB89C63589074517A6AAB1971ADC0482AA337C1439BF1E037AFE9D2F0EE3808A2F957A40FE03B814CD0443826F7D0246CABE59557D09578EF9C68135FC7BF41BA0C1AACAEF4E7BB779D627EFCD241EF0E4DEE1D66B476285FC539C7958CB51B3399549989588A171DE4769DD1786CB7C8EC157DD5F519D6FA3A735DC1E300776C883B520E04874EDF3CF61534A43ACE7DDB580C7EEE3C260E088486A272E09877B34B67B4840380DC25E67F405043972FA27CAD27DECFFC176A62F8B477A265AAEE6E47A2F073605E976281D14EB6C4468A5C0B568189CC2A6251B68ED8F1517B620E88B346CDC778143129F97681C5F658EBA4B8E6B75E7E3C484E96C6C93F47C5D6BE6DCAF1038BAE2BE2172237967B62CCBE229BC8C982406FBBA43486C60FAA200CCF95FFC3A51FE71CBB74D9EAFD6B3D1B4EF86FDEE2D2BEC70D58C7B0B7319A8E2D834DAD12FDDCAF9E2D8F69CC5E82A38B03C8DF9750BBAB3409D274F677402CFF1F33EC9073A1EDED464EDC715EBD024B4BD11BC5EEDAB5B01E74A6D325D41D781696792FE7AC6B519DC5F84F050A43485415CE0C71CB99A556BE376A977E66E68A136B98914A790A2E65B40B3CDE63479AC98132631E2F9452EB8C4DD0D84AF5743791DC80E7F64CE943C1DABABB6F47629B116CABCD4F5E9B922B1418657CADF0E2E436A63B6B5CFFA1AC3FFA1E67106E39B5B689A30C4CCACAB50819296F4FEBBF70C2987090F4BBF5AB078AE88350A4C3865A75ECFAB946A0EFC84F7F27410FB88B4FA6196A007919EB47724BCDA59A484968686C3B8B5DD66F7CFBF599DFD25945EACB8060BD63B73899F7346850D00E530BF2816454A8EDD52CB0E4BB4DDE31F3883CB597F748CC9B6C5BD7C24E2BAD857B43B18BB4D4C5AEA2FA0D99F0FF878B787A77A6B6FA3124F9FA2F67199FBD0D4D3EB7BF41984DD15F94892B57A671B2649510289583E06C817C4910C5658331C9609EA5CCBBF2160FAD73F9497A0C9F7DF28B7A236E9160DCDEBD90209CCDB'
		},
		SiggenCaseItem{
			tcid:      4
			deferred:  false
			sk:        'EE620C920C1B1DA74DD53ABC96E69B2F3E7637077F85D7B9CB0395D9FF69EC8F0BB877F569B56162B9DF9A6A621A81A6AC441F7D3F642116EEB752A9F823723A'
			pk:        '0BB877F569B56162B9DF9A6A621A81A6AC441F7D3F642116EEB752A9F823723A'
			message:   '367774B2E217EF33D8D42EAE3B69EB09060DF42FCB408BEFC787C18F1834CF7873EC07AEB460CAE73EFE8C8FC0FA39A7689819F5E182833E252912ADFF2D326563EFA9751053A11F02D5B24F7EB118DA34C1BC4A9932671C6118015680CDBDF04E0B41D9D56E6925E2B328499FE5562780927ABD1D8070A4C87EE3797884D32A1F5135D4D9996DAE7EDACA0AD7309A45927ADB53F8DD4183E01A72421DE700ADBEFF79392AE8A25BE6729A5F0450BF3BC1006178319129988B60BD7CF45321183ACE5B966B5C45F3F30CE42175CCE39D9767963E003A7C1995E59670DC9668CA94102CE8EE56A2573F62B3ADAABF7E21D09A125D1EB62966B64AEC0DB38555A6BA8FE1F4EDB437AAC4B4F529A0326382F349F5323C235976041A9C2600660B348C54E00E41716BC6CC4F80772C2D805370ED74BFB9E1FA9B9E2265597A04F9442C21572186D46F6709AF1437BEF7996A73172BFAAA3756E37567E3B1D87475E1873F6FC598F36A9BE71EF710C5700281D43ECDF0E580839BE7EF15F170578600BFDAA7C1796DA84007107A2ED33DD38A5853085F7535BB2F00E932403472AC624DCA4E99FB5BD5DC9D4225A0AF84841A3049641CB9D3CB0E73A21D4E4946832DB12AB2585803D4BC70C13240432ED21E377C87B79F5D8D0023A69DCF18459ED08369CF81A3BC97B701047A46D3EEB410723593E816069680AC5615EFBBD6C0EA08062FF83E4454CB659EBE36DD3956389559A5D930A6D6B2620DC6F788FC56C03A588029274A69180FC48EEDB9F98E734D9DEB1196FB43882F5743A85D638FF38B772F6BACA3D5816A3CD4732E0609A5B5245B17F0E1376AC42DCDFCCCD454E437BDF3C39E4397A8B4DBF3CE6607B5FD53107CB247C6B17E3BCEAF444C8A5D5E0A3B7AE4035DB532D6A2DEA1607339747119862A325F1FB1A1F62154766D4B937D5341A07B2616DA3AAF11677853755C2325B1971DDBB14CDBF60A1A38F0E1E70957F4D5D05D9A23B1A405E4ABFBA7AC115945575555EA722811FD154AC77E3F93BC6220FF86B6687D07EC074DDA5ED90B54E2B72F75A46C77F45C87C6172A9DAB53BF09D4B301F31174CCFAC161668598C42D74652A9352C637D3007AC8DD4A01AD68B45FF79D38C947E1C3C76BA34BF5D64FA4612C4B14081E0072ECCA3BF337946564AC5B5BE8688EA1B13E9B71C6A9BFCBB5BB15DE66121510BBDF05C76AF8205E39324C0BC08B0AB93F935E2919D9DF78B335331396CD97B1B71CE6F221CE340F68B44BA6217301E8CEABABFEC4CD2DA1D127969E08891384D86E7EC274D965EB9122F7467BB1A049D43C9CA9526F2036DE5ACB87BAC5325FFBC757C1BDD5256B55FE6EE4030CFC9DAF50643AE80E4B30303B979945BBEAFF06FB53784E4F9A397685B89EA0507176F41042A4C5395A4E3FA510570F9BF10D9C0E347583F0AEF1F52A73435D8BD64192A73436C8860E3B70D668FC409063E9C915297691041D28470B2BD474CB25A8A251E77385BA22C684C67AA119F5FC21FEE80F823478937A1AB9F1EB4D9202EB7782F13DB162D2D8975DEE247F38E238F6796776B79D2A938F98D55793BA2473EBFAD9FB2DF39A655FC61F5E0C2213EF1184A67106EDE5517E1E314CC8319FB7BCFA479228F3BC9DEA6D649CEEA9B2C1E59E883372E16D328C01EFEA9185D2C3630D08BEE4F88E99B71852731F72526E09C3D19BF403C5C4B92B8AB68D74B63DE1830F4017BB84B6397D3637A5275E17B77D5F47C2B447734E1F7A68AEC717EE50F89B7D8A09EB680A944F3C7613E43494397EA46306367C01994A03238F4A89B9AD4B8A5CF2513522C24EF830490C98229EF7F951D09C9B82F770DB3F0E2A598D808583AC06D28C32CF75FFA2B974727489114EE8D7093E30F7902F7E840498C2F1B2A5BB812233ECE0D15A0FCC931327EF5F44A6ED4A3F254105CF3ABF6C042985CC36CC9B61D4CEB83B33172F7F35C6CBEEEB882E1D8F287F411C56F1EC2814E8898F025ADF15DAE873C47C73BE675D5BC026E881ECB314CF91ACB13BBC417CB7A6D596DD9187F1D66C74E2325EB92BF258133368E0BBBD206D93E1D1EC475D56F6DA2CE95AB66EF38EC83CAAD48263727D9E8219987292D3BEF094FF7A809FA81EB7B4C12CA891DB2DCBDB728E7C1001935C528BEF7B0DAB9C5891EB929BBE6A3BCA26E584F6CFCF297295A51E2F2C50DB269B39EADA73459C38B8FB77BA4EC371F9A2BACDEC282F953C6562C1A9E3555409A5E05F2F63DD85F3D1AC26640C8FD5574F0184805A8107FB694EB7F8386DE5DF60844A231AC0FA263B276D302AFE8B1C5AFA17C934B48DF00479EF5E03C01A3FDD516397AC305166CBB935E8710B7459ACBBB853ADC230C31BF6536B26C6E0700FDF3B9F5737D8134DC48C6578A9E757E51624E4312A1F19F0BBCF84439E2A571EAD9158635A6FD09FEA7DCCDB207FEB7B970A501DFE1EA1389FF9C70877FECB906785F79462EFF06641E250CB57B8E982D7FC416ABABFA4A526BB524AD512823A4924940A01C377D9750BDCA2C4C7F4F2439C1BF93814B4FC90F957DAC865721E8514924BAA2D1FF3F67A7F6FBB349E7D961BAF4731074FDB703F3821B66E54F47A98D762458A0DF3E44C0188F0243BC81A0E481D5AECB65D76D7D5B8200440F8027094F7FDB88BDE380934E864C5B346F85825F66657640F8FD41AD16946FC1934664DA46A33213F04AF74BEFC463191A83FFF1D1E755E5014FF2B1EF7908EADC8312E96575C85F776436BC5A8790EBBF31261F7F4C54B63FDA401EF2B978270751C380A0125A30A36F3E369D85CF515EF56B67A0003CA013C30BBFA67BBEB59AC44229D8FFD11A98D62FABEC68794B99F68AB16F12FB497BAC70813CE306C31B2AAF06D16957E9A6DA7AAB59A84C944448A2BD3EC9D039CB138330D987F51371795428FCBD844CB3C98B4F4CC66CFEDD5A0931F6783C6F439BC455A60BA33229C761B69719EE5D7AA9357B3923D59F79293C8CBA1EDAD32FFB42EB1AFEE5E934C4632255D62819E6C340D15B6C6A9686DF549BF4E7F69CE9C79CCF33C520CB8A90E7A3BA5C6EDDB53164A0BBC4AABCBA76B03BCA608A1C682D8EC4B3ED5B5B740CA5F629150D371B2F0C8F045EBA788C40AC8F1094C8209700B8B79379FCC1B0790F663D270D5705D0C08291112D20E5224EA0AF1BC47362D32D267C0317DBA19D90217F9F9ACAE14B9AE5083B03C42734CAAB55AE5F50AA7F05D7F1EEA290B5D8BD94D54455AFDDA44EFE7C6EF268BB2F152EA3DDB46F227575D54F687F304A0753FAA3BEE33C536E890A0D81D610444530612EECA819C35143C880B91E56BE5C70428F36BDEB90341B4BE777C0764DF68E5DBF2D8CCA59E331519A73606EBA6081CDF82416D292FF8EABB6F1FD04B2EE4BF127C8C7301A7866A61940DB1EDFC24DE47C735489F7A616765DA732C0894AA275924020F8550E314CAE0E78B975EC42E9B2864F5563DE3158B11C4E5BB514B4820A410B22ABF06ACBC8B86828FED792ABF2F7D54DDCACC6AD72DCF8CFDA0A0506377781088845D187C42C022A8BB425A9DC1855CA1AFC099B5993688D883EE7CAE2E3ED24816EB458B1E039D6481030EB5A80FEC1D4E7EA249C12774C9E9377FDF24A4ABC9F803ACADA2AB2051095ADC0E00711002CEA152DA07CA4BC399E8373F54A6BF5E120E27B812BABEA158A9130CEB0EB12076D386E302BED71FBBBE68614C78FA1C67C71CB19187D655845498DEE90782024983B84EC326252EC0B940E81043F6F188FC146D10FBA42E224A0A28ED97D8FBA778A4426A82197C352CAD36B6F99F8F7D8576C1032A7AEEC622D1DDA35B5B6DEFF6E1B0D27376FEBE17978BE96B51F428AD834804C7F2892876B6E081D793CDB896A107EDC83C00CE7A88F5B3A3647D0253B53628130391FECF780E734579470D4B2E4DE85447DDE4AC5C0858F158A1852A25FB1EA018E6E4895B35A520AC2B83E1E70B44EAA7284ED4D741FAE81B5A051D2F2070FC28F45773388F7D96B1BBED57F0734B5DBEB44A96F847956F5A1C19D8CC56DC9A8373553269039EF1BF471B6CB155043433D1730CBBF3707E26C076D6813CDDCC289FADF4A87E2F32C1068A68C5BC30D1F39A15AA2305393068FDB0983560F84AAFE128E126F7CE487B9711F524D87BD759AC3779868DAE5181D3EC77C7AAC9D2FBAF4041938A7D2A149C37D156BA0454747743FF32F4F9F022BC6CA422E3E4B26967B0282CF04F9CAB696D807DD10EED780E5AAB5D323AACD86D31E3262993821CB4A264A87C63CE23A0326CA0D15D54A092CDB66501670CCC58A590BE733DDED50E51DA25AE8045C5BFADC43F06047DFDF056630769906E8FC81328C2288ED0647172A54F5B45F7F6D520F56FF6D4DF8068B94C44A14F48B3A0356AA5761BE5B51CBA13E685E6B73D9B0557B2440EC433B89EDD0E43ED1F85592A35128292FC2CD33A7EBA08981F46C79031C0D5A2DED647ED377347B8EF9A751C7EA42C7ECDCCC62C5522E40C21F01225C7328794A1D8CF6190505EC358285C63C72989316B8EC2B955767AAD37D83D9637A0E04BFD3C4508D6970D90851BA3CFCF1CE55F8749C6A77E85D1E7E0A5F99EE1E4DFFBF72C7FAD88107B3236413E265E5B5230771F7A169CD8787CEACE1851CA44D2C342012A224C5D7E015F6280F602BBB6F9F7C3E3B3A721FD224ECC0A0612DB95B63840E1145449F35AD2223799FAC649F4D52B2C5FFB0A0423167F6C40B8502497FC7ABD4BAF8B242422DEBDAC4513A1BA0CC25736739131F68C90A0796D163990CF7DAD9C8156B72C61A0F02C0090B4B6F8D956F1E0F314AA163FA166B786C4130BBE3DF9C99A9463B4372A883C48352DF757003229454E0C76773616B96B648B282D7536BEAC0EF80C80372FFF8B214D555BD21C12EC4080F5FBA5D793A0E3EB6729135D958B89CA74121E69C544081C4EC9B69D57CBB53B8A0AC24776820B2AEAFC7307A770160CF929E8C828CB8AB7431B599ECBCEE8DB31BBCDAB9882F35CDA463550FB4B37A868816B3FA7E7F658B55ACA69DEE6711F4D6F53DF187E8E65698FAF1E2340110D8538853CED364B849AE62A26E75DEB8A6559910D59BDE1EDBE5975F26B913EE080B1C7CA70D678DF7DAC9CF96C4CBEDF811AB0622192BF4C02F5126615C83137E09673A53C6DA515BCB2A0190AE4E2D0BF8BBB9DC81F77F357033815EC34911DC6A7DE4F1D7D6A3CB87982988617503B0AFF9AA7E5F8DEBEE59023A7AA5D8E3E4B26315A1FEDCF5A32A095A7DD5D847BAAE2727B73DD43F701FD3CECD79DDD4D205FF60A92FB1D7D7A0D8529EFE0BB227DFA4488ABAF9E4130C4553C6B4A67B8CA8587997F0176EF6B1E2A111F74BB573AA7363F55A8D3A7F9760B09EA899BA41FA49EAB37F6CAB43A9A317E5697B73CCD40C606EE865C6831BF8F4AB5B08A9C9C81A9D7B1899800AE25C6B111046689C0C1B975253825C87B4F35D0F678D9004C4282BD2178FD87B5EB3F144FD7B8668F86C28FB1D6DE1F3ECA4FAF104DEBED3A1589C96AF61083506A4C03576493CAFE451DE2661415D60BEDB431FB4EF101EF9679E2A2B7ABAD6829A4C6ADEA0CF2FC4AFD024FDB84B4F72B8016A479ACF431F9EE64578F15FB476DBDEBC90D018C0358AAA74223FADDFBD072B7B3F31A26146DD4AE77104AA7F23F254AB87F8569E3340ABE9FC06106A76574A237083B6DB7766A4E77E4C00D164A68A429A2436F72A9BFEE60D29C7FBB4C93371E61F25AE34EECFBEFF813A2226B913C3F1D523B9D920329621FBCA3725A468A87E378A887A7C17CDDE00276D2220E1D760FD902D61B1B96097902A5CBCADCF26FE6C53188074B19202957B8290DA365C5876E4E4DB5704D1401AFD3C1E1A535992B847688D3A4E45E26B847693098B84DC48770FF751EF35C4D042CEBAA40D870C0E9C1C6F02A4DF76DC46BA9CD9B192D9A7D02BA16F582ED4B66B2209C52229261140449C653CAC64286F5F80B3EC20025C93DCCD23985C433871ABAF08F7E62BD76E78F9B3EF6D84AD4F39CBAB5756521A3AF1AB5E00949A4A088BC2C149B3622AFAE80A4E4A3D5E3F2ADDB822A65BB4446CF8BC5A1126BF78B733F14DACBF7B076C61F71B9ABF02F75BCC74B01D518DF9D97F70C4BACE9CF1F3A4FD4D24AA0BAF8DC58434558DC3DDBD7728BE18B32DB48115E7B85F08DCE0964CA96E9CC06E747A9D733B061F1FB127DFCD97BF334E9D039A1D931E763CF1008A43754EFBBD8B1ED7E15750314EAEB9062E9C09ED7AD9C1E85A4A5B8D5C5BE4C36C54BDD8B7566BD7753A0D00856DD469106AD221C47CEEF14E065229529411FE57D59F2307D96100CDCE5A59DB0FFEAC63AE116E4A4CA8FB77C5A228672995CF93E800740A481731D92C7E6D6856C6E02EB952F853A5D66859996B2F0B3A2D3C2BB2B091F01D55B6A6751420B4F294E2E4BD628465C1824489F091600EBDA6ED4D23500D49ABAD913DB8B9E5FA6068FB0979DCB2277A5F8BC00A4D9DBE936F505B1E911DED9E5CB16F8A0EB54D425EC79E4FF37E1DF1FBDE314DABA66D0D1B4C7E07284937F73AFCE7EAB4135890D96BA0AAAAC9DFED678357C905289B34AC13AD575626BDFF723919D35B758553A7467636EB1920C893C42DE648AA2054D033603976FFE74FA28BB3CB9273A18569A063357D6B781C4D14473D66508B25F4AC46FCFAEEF40A7BF3A253256DDCEB019436C3D0150117306B186AFA634344EEE9397F5EB3299064335A8E82A877657F4190B9956A1F2E2B95B0248F584DC672250B9CD35C3CA24DDC2DEF432CBCE08F97C34829B569EA760CDB8B55677C82229DAB3F98F6FD4289CA6F0F44853AF721158BFBEA60641D549493D0AEC67CBCDB72747E13DDF60B93ADA89DD2CE7F19DD7A41D22447F4971BBF0D9F0290E0325841CDC39F086162E7A043EEF77FDC622396619EF8C4FEA93603768540EDBBD79CA00DBF30A2A03F094AA712F13AAA92345E7CCE688CE266010E664F476ABD8EC33519A20210C09064DA1BEB3AFFA79C52CDEFFE6C8F1CA6521FDFF13315191535D21298C70D50245CD94D85333485D0FF9964508FE350E5DDD0AF62451D79A25F4F2FB0D09735B71E7FE1CD64EA86F172250EBCC768545592F33FFCB46E943EA6B26FBA3607F5FE562BB8E438F3D90DDD63C0E94C2064CF0955B8D6958BD2C7542AB14DF85455430E5ADD2C275DAB5BC9D5789735E8596800581E8B4B04592347E031E44FA2E3560AF6D1A588651717E103DAFEBF2AB7960F00F0DBAA5049EFF055914E758C5FA4C437C1ED8E68690133C8EB84E45988E92EB770AF57A78DCCE4500DE1764AE0CC98CF483803D64D8FA05883382D2E300E4707995658F8741C6FD5C3CBE80959B6F118B32457CFE0C80DD997CBB3FDA2A81BF5FAC001D1E55BE3A007F4AE4B5938143725CFD65BF441D79B384E4467BC77DA621741417DFE26D899805C11B8533617DC2370657D1A33374C3DFFF8CDE573FC19BCF181711447A79B3CE08F3B8E058B210C29DBB891876398B265C5A5B2157A0F979FCDEE6713F60F2906F47DCBF9A1F395BAE35F7393B98ADFF8951A56D092315E5B35200910DBEF794F4C4B02439147701C764456D86ADCCFC70F42F37F5E654206B16D4112000BFF3A37DE607941EF3B8889A535E4481FB88642192CDB19B12DBCC45422CCDFF9B1AC38AEF8235301E02C2E1D207C12166AD43A211BC1B837D92001C38B320B69A5BA2157FAA2E3E2B75DDAD512F2D12F704F862E3685B3D3042351DC161A6FBB01311001AB9255F10260B6CF94BC6B2B0C17DDEAED0C9AB5BBCCEA40A3F6536E1D7F917E2DDD475E2A733AD14B6FAFEE73F5D269787D3A92AF3DEEE2E070743D31F23F44AADF20DE71565827AF49F3AABFCAC1182385604CB44C4D4EBBB8A4829AEA1B4F1A6FB9451E05FED8C9EEEEFC8C9AAB95031F275D3149A464143ED4603F22069E4680456B6FD4375AD2918658B0618D9028E3A4A17861CF5FCB29194550C17A50379F6E1A2AC478B7B0AFBF00996F8D3D843531A9724E2DB4AA603FD88BE7FA91922FC83DAF11C55A9D26EFA61669CFFB01953D4B630C700FDD0D2BF02F05DEA045D56A596A8ED2B17094B5E24E0AC1C6605EEE6A9830670C7932CC71C335FF43193DA0D8302059EFFFC58BCA18E932A98EFF361E58E7EDF6AD9A79C47EC2870C6ECEDB80A440B5967D475276371496F2F74B445A425E11F4CE5518E5B6D727424BB2DEAFDC39E4C349787C7AECAC4BC680309BA614D2CF3D7EB7BA89040F0EE9B23F2272DB272382E1592D018B90AC78DE2CF4C5C0E9716E35B9C70FCCD61C768A080B892529E384F65C8F9640F4E745B7776F208588F1BDB8479CCEAC19EF70FF7E0672D663F04D4D8A4EB2A739B5D2787319AC571BE4807AE1FD2567310F350F26DFF6D76FB8D123B63C7A197CAFB56D03FFAB4EEEA7DF64DDE29F35240379F4582F46FF22D6782E689AFEEB596E5D8132496AAAF39D2E7DCF19BDE7E739CEA517C377CA20E7B67EAAAEEC1D159E8E8BCA867EE2B891C7DFF967E6D95512DD44B81489E7EA2807A13C134CCB7D27E5B5F3030AB48E76C991BB61F22898E291E77A5944FB54719EC54AFD5972337331EB908FCBE70A47ADFD0FDE5988ED42AE9585703EAF037635BEFA050C3C63C97004EADF6B47782757B90848718A3088CA4729CD3BA3881CBB0BC7440E61F0A64571688A01A789D852C123C6CBBE720CF2F8670CE2A94AD89EEC76F52FDAE87B7FC406E397238131541C76868C170931F0E71EF6ED707A4C64FFBD82D8DDE4D947AFEDD4F072F411FF447D5CF5BFD84C7F5FD304B4302B5DA8F7668B357075C1697C3664637891D3FBD33708DE1343DB7AF2F35EAF5E558E04515D8256EFE5265D4B70398B434F62BE826309CE3FAEF689BD6B2A96D31CE9A5B1A7B2EB40565EECF5487D09CD88E62D9A21CC37FB4FBC0448C2BD4ED21BA5C889F704396D0CE05EAB050DFBB33F4C6ABA0CA278E563ACC5E11FF820A509F1F344304919F3902A4CAAB1ABA805AD2430F35248C40EE9F8C30107C997498B0046BD0398D7604FCCF2C0B152EE36BDCDAAB731BBB540AF06DD07B959B092FAFDFDAFE265D347DB62AF17996305C7008C6AC86C823788A03912E6E0B2D2FED49C33C719FEB32896073979345589B1EDCDCA8C58952F2EB5179EA58E695F14DBE37D1324F384CB08B36D8BB0FCA04EDE91504FC7BED241AF68BAAEC9CBDBF392EA65D49468533E1D823B2AE6DE877FC658615A5CF20F41B8117B8821925D43EE445A386C66974FFBAD41D6F09A532AE0EC41170FBA37FD22C23B3BA85EEB5F593BB549F9785C077F711494EF3213F34D23D71CE1B67F939E53B0C87E16B110422109048DA04EC7F932DD8F5DD640E38AB942696F3D70623042FA4830554A4CF0727B3015AEAC9F8D464A6218BFE688ABF11DB863B192BD611EA33A4FDC0E43A4F63F345EFCD4A861A'
			context:   '03079F62E1B44E2AC1CD205468B776B6E1FF9033A021C73893A8B65AA708EAC07D4C2F9422F808F68B0AF481F2BD4075FEC557C14620DA329BC25BEAAADA35B64E1311A92D747C38C1D7537A5362FAEF936135DCBF39D38FF55C099E31CACEDE8548E4EDACD3D633A216FB1AB0CF8EA4618CB478B8BAFF3300BE7C03A81E4FBCF1034AE2075C7B47DAEE97BE6CD44D7260B1BD8086BFE2CF2AEB4A281BB02139D567EFFD42EE561E0D3B389B89291F4AE697B4C9572423E0018CD05D7A8883128920E88B1F340A147A15A5AAA0E45BFB49C4B19EC3AB5ABDF30E324C03D133B2E5D87FE525680F97'
			hashalg:   'none'
			signature: '8D616B954C513D1979FB5C4DEC591DDFF8AFB34190170088213890085547A5926EDE1B37B055E342CB86F378F7AB9011826ED877FB73A68F9E7B88B52AFB5A80F82011506569CDDBBB451E9DCD94CD4A3B4E377D58BB95FD50B852A24B98DF15E1F1655A16460330FA69B7A7BDCBCAB31AFE712062B1D7F14E8FABB406953CA137EBE9C0327ACD67E2E25A5D9F5486344BDC7709FB37B9674932B5714FFE55F64176DBA3D23E92EB71EC50F2DC51BACEDAC816C3D91C4DDC71FC6DF9FDAE943173B632EC67F91CE7897DACDA0DDC4618915E23CA67C07F956967480444F7C40ABBC5F56520B981BF2B89C9E437F220D8609D4FE1A0D9EF81296F0D877B47E7B4F3B793145B4373755C8EDC971404B52FB28F6C4BF9D40ACB565F8BA635A562FD32C80A011BE6A2C13E59279D626EC82A57E6C292E5E739FB2BD85245433732C60DDC0A14614C32CA36DC0F7AC516B8061F286F606D9C55240381B7164BB8D8BDAF453409A45560D90C8821552FE43826FB010C7CA7A9224DEAD7990A9F5E41F6E47F8B2E7296B005B9B6FE4A8F89E2720972423AC2D5A701ECB2002CA21FC149179980C89DD5B04B5D8E970FCA145E4821F3F052C402C341AAC80B2B114A49D1AE29E62029AF4D86C62C3574669F2B04C399218ED10A3A34EFDEA5056AAA5DB7D6B36F9F9D46B61D905F9EA62E6E50D34DA06047878714A6D51DD3E2D33FBC0B7114188D29CAAA49198A69CFB39F8D65C912402825C573363D76CC1C4F467D92FA6EEC070E8B88687D62712A2B1F6E27A6D787DDB9B489FD3BEBAE8C32E6CA1B736FC017BF7F31084CFE85D389F4124CF23AD3406E165516F7822F34B263D0FCD0C6E6E265C678DB3D1CE7F8DC242BB24F9FFB9815DFAFCA9112F4138716B3E88147DE1DA63393EE3FFAC8493AE1ED96EE4B0D069FC41405D57ECFC6BC3412F5257F887B3C3A0058AF0FF4795FB4CC213DDA06B0ED27CA925EE4C6238F89011C627EE40D52B10E227A75CAAA259F7D0ADA7F5C63D5CE9F4A8F2056680B4B77401D5E721AD581A5EADC44A8D73E2072857692092F85B994A491D4D977A2C7F8EFC4C5005CEBC58617DB811BB5FE49D16BFD1EEAF0EE9A4624A64D76A26A8DBE8149E44EE84C185060BF80626270CECA3450513A9A9E476D612159AE5A031247F58D087F72387FBCDF62DC546110F8E0A521076636062B6A91B11152CBD688C7F5ED0FA6D99E0354974F6D39B7D294282BF55B878914A4949B7703EB1D98093516553C4F1E9479EB71F932572462C625B04E2CCCE2F9C7818883989D33C427C1F36964498E2313A828F875074D6B06E43CB50DE40E2A75B7363C5207FAB66A66593512626F336A1CEECCB273A190DB804499516CF938642F6C39A4A632FDDF8A78E5634505CF2486EA611731BDB4284BFD9238DA8D057572F4FC315F9944D588FC18E327E54589D62BFC12989A8FFF9F66A2BC4F5FC8CE3EE46406D4AD5EE9C8D84700517157F49613B2B755C5077CDC73C8539E1DE3D7EEC0DDAA2437B483C3B8ADCECB1A55D3B03BFC7DC5EB3C7785A153D484D83594A1B7CB4513C83CF54306458F4BB8B5572219F39C090DEA82FD8F2905EB0170CF68944201A05BBCF978017728A3AF607398D6A8A88CA4ACB717E7BF039C5A5D34DF8CE9B92AD694B008E7D645CA6CB6060C4C0AD2D1C9338A38B5E0CA863BEAB1E60981B189B28A2FFC5CD7D039929882556B42C74D8ACEB2C65684BEBFD1A35FBD3D9294BAE33D56D13EAFAA60AC4664C3F8B4A7D2151DCFA201DA79655A4EED9EEAD8E917579EC68C4CE410CACE1E615EDB98725F93FAA2EA8E82ED95090776C09C9912B1C48050B29DCA99CC0780EC26204D6E1971CB8A65925C30BA47907A9CA1D32AF9FA4EC1A399F4D9D80C8F708CBC5A9F4548A971CCD2ED670B842A8EB8DED8B45D08E6C648E918D3BF6E8076F2765456FCCC610665CB3892BAE6A891A4F74FE77BBB86B48F122359F695247F9B0C5E07F6DB82C037F3B8B90BEDFF39381CD4CD0592E3F1CC9DB754AD5B422686449D8E1700D839C8634C805375453406A027C7BB6DDBD8A201FB254DC2FED6E70FF19EB02AD367B99B5DEB7B37BC1632531509EFF6599508B33EBC9C03096E782F921E0F695FECE9D21B24C7231976C5DC65A4702036A0E2D93BBA1AEAFA7097B03F7C5E52F053FC2261EDAA2613CE8DF7D46D520279C06153C2566E8D248091823DD068A9965127CE00D1191ACA5C2CFAEC2478EAAF7B601A89A05E8CEB76E24E42A23CDDBF983A521C60E827D438A363514A4FB3B3CCF9EE080C515360F124215CC40C2579B598ACB122C11AD5CD7EFF0F493A7BA8CC3C294701296AE914BD11AAFB8F77E8FDF0E2B49BAE092E9DE02B78DCE692E8F9A6AC8FDCFEE29DD8A844F9D989A86948DB30BA0215B8BF5C6DD915E9CB91288088F3CBED297C18EFD4F21F3859765FEA4EA31E905519B1364FAFE948C1F9458CBFE02846D36096763AB3AD79970C341F5A8698790222B00A87BEA3564ED33E9163C19A99D2ACDD25C62A7E459D02977AD937CDD69935705DB49210D9C0C055FF58E9BCBA082DD041261F3897AA72EA52829A283B947E3580825BCEDF7D313C104AE29ABEAC14EFB7012185A67B152CA378265C23C757E402EA4358F527AEF2D1557F27BB0864A30AF48787C246F16BA2248D0CA3F7147B3AF9EB6C4A9E5E65D05D86F6F1F40D8321DCDEA86F2E5CADE913C9A04C5DAF1932812700C900F74628CE263BC1ECB3FF375E6F8B95E4A8C714FC267995B98B09342A1293FBAFF4D140337759DA3F774955DFFF2769CA54E58E754DAC8C3E1F6584275B1D3F23B5C59392E2D7F0EB0DD7488F177961D35C7A8B309DBEBBDD54D97DE3DBFF02DE7DE098931B144505C0F1B907429C83EB20ED791CE575C8C34F9439F5025FA29F5D2A6F8CE0DD5A20FB882E868B543BDD69DB556719DF7574BA6B2C72D924C8760B890C5309DBA90218141C6870EAB9BC814997E4549FAE66D920FDF5CE98F4068A337EE962A49C89B0FF75BBA27E5C8FD9AD4F56D7D76E94445F5299DD1AC6900F4252978CEDC6DBBC412D97274DD7D10798CD7B3A5291934DA041D3C7943440BE89103339B0A6DDF4C09943B0D99F5F7CD77B530873F2260206077DA2FD6D6FDC63195B396BCADB93205BB4702DDF0BCA8B3D839D16E33078E5BD07FA38418373F4C6CE3D73B596DE7E7712053614635F02C9F58A78651065C7D12C3530339C216E1C2802F223CB46953A886D3B04A502EF4D0273C21E3293923EDACA6431A29CFCC050F17D79CB959EB1E37C7CDA1B5EDA67E77A7F461C653597FC99B7CD5806D7AF4AC1F2AF074A93C93D88ED4992857E5F546983C09DAC2637928906C0E6531DC443B62CF9B8B5A19A3F9F9395DC31060BF65FB9A74827D72E8F9D538E551F47B21890823663893626AEBCA98DA031D3036A4B1CC8D63374968A52068F75E6C73AD7C6786C215286F1270510EEE6B48D6F13AA7E8BDC36DEFE7E36BD5441188D87E10A8F464E4E190292EFFB7D62E405EA669AA98907065995B8A99CBF4A363BB43F7C17AD57CE15388DDF31E630414E1257B8AFD14D3ED305E9E74F948BD0603EE298C83AAB985EB91A8A2E05E564EFD9FD114E0E48E144F54F7C2D9B2A426E32935A2D84D1FEAEEC78AFD8A6C0E0CD6EB043F508ABD8378A9EB447F1E77744828DE304C23D249A5F1DF7A70BDA45F7249969262AC5AD37B771B983A496D9AAA65DBE3D2DAA8D4579E849D835AB6BF758BE3E8D1CCF62438D97340913A44DFB2719D2800B842769DE7810BCD87AE6E1351CB79713B5DE2DDB9C40BA7589533A9EC0F9BD322BEDE26361EF3CB0D6A21DC0B41E0AAEC7CAC0EF68F84252F6D7716993F1CA481F8778A1C74B5E07005AC3E6A08A30A3B4607D0639C781EEF2C2193C1777C556FE5B3DB98134D9D07390293D2254F242974F13D41382CC4F1FA1552113C27A285A127547F06804210E2FF3E102BE903A96227FEB2C6D131A61AAA217A3EA903018915BFC90E50F5076E34A20295190D18C1C0E5BEE32821F19347645C97B1626643B2EBDEE7980B0CC7B9BD859140D5627FD2E1F3A5E07B422C10B7701BA2EC208C186178CEB4E963DC68737B67A5B75F7B8B0A01F4FEFE73DAF8ACA044BE30C6017B8217A53D05EF66348BBF4398C44C37E93910D3352A90E390456F29423EB1D83403DF255E3186D9893A67DA10C3D5F5792663558A843FBE12F12A51B57612EEAFBE56F2113A231716AB99B2FB16E0B035EE68384E29C2AAF3F710046037A6FD90B71F906AE644FBCEBD0D83E37C90D404855BB4273ED7E62870ADDC0D7F84428D71410EC525975BC2106FC77E12C9684012929E3D805E3DB49074A2D768F7480C3758CBD23444BFFBBBC9337AED6D9F5099334F235393CE9DB4EEB8ABBADE4D6770BDCDE3F49C502BCF84A942538D9ABFE4F0981953BA4BABBAFC78C4692C928D4FB41413E12CE5DEF23146C6DEEB28A87DA83E3619EECC403040EB75EF38861A4D835F63463D8530B679EE6A8906D9AAE1F5535094DDB86D6B5E1883140D5A65B143D5485A4B60637AD0F0A1D1CF38B49A7501613BF0CD9955191E0CE704DDF014AB7C9466A32053E70F074D46EB2F6AD6E7BA2086D39E52D98C05862D79018B55DB8F4E2BBBC485F30FDED502E3AF0616C39A58D9B680527642BA6605B164CDA02782F16CCAB2335A3FF5F7FA7F33EB0EF0115832FF93BE469A945D72BE7E029ACE425F0E23EF1B0EB47C39415C813869E6505FAD22FDF6B3CE200919A40CE19741FB4A71934C61E537DEBDB0C2795801DF5247D13648B192E4A2D3A6AC43378CBF59621FC0C2E4A17EC1003428751D2EE10B530481B5B6EFEE5D8B2757A9F0AA60E6C4E709454AE6DC81432EF673A2E79D8E726CBE00CB0D291D1FE4227B0D393382A3013334608D65B8172DD6C0BB2594C731FDBCDF31B93320E53BA494E0A2003A4D27D723CF2A8945D204B2EE0B29A12348D511A7FE81C43D8395E0D5BE9521A851B2872711C0628810F8A951B42CFDD89B20CE4B3CFBADDFF5A0DB96D9AA9B6E821500CBD141436C0C2BCFD1891C35DDD6F74D7CF350E04B63735679612F59E4A594C164075EAD9082BDCA4736FE230D6C9DBDBB2DD0426F844DEAEF20E8261A4B2E0DE72146F0506A582C05CB7837D25BCFD23877F3EAAF220106616E8E91AE73C401A3C7080E8DA0484898A2D8709BA276DFE97D2C58F09A20A59D54C4A75E4E1EC322F7AB7C5842CE42F21A73CCFC9853FE69DED74894EC0719BD893B6A824A624018C33DA604E321D61D9C44BA842776E3258D27A3C477257E73119370236306CF18F2E1473D6E1536524FC4C83E6F8E93444FE5EF68E5A9A7F048111A4990F0A2A8B3A9B5EF5D1457130D541DAF9695314745A9930B19627B65AD7C17024175BE0CEC3A64FFA344478BF8091F370F1C6320D0EB8455E24938A5E91633F60A842E7FE7E5A907B22D8686E1999482A474DF91502363EF0FFB11ED8B2CFA2A8C225B156F3BFFC117DDB248DE03A1C0E4898413142DEE1A40437980C21A39018524C8FB5A378BBE10C14DE73CA94D7EF03BD8B9130A5E6C105675AE86A8579F0966ACEC7F220E59EB5BB30FA7F5FBFBC44F848AE9B0376CA7AF0CA61F270533E12BA288E71706F14FDBFE8978D282C60D3547682C01B759919C712B54DCC99D901F60D63C9933BF0E52D25CECFF663A61EB452B4017B20BCDD46202CAD87739DB6A2FF0017201F4BF355381087997FF419DD168A2D70F9CA95ECF59F6D58E09994072B0AA8A89A2C899100AAE45DC70B8C0B33CB7F7247FC40502E4DF01B69785EFB7112EA46B8307D3BBEADE25F752C7F631E16FA7F3D9DD218A840B477CE51B943D5358D9981C5076105C4190EF830BA628B7C4EBB98D27AB5753D4012537E21CCFE112B8F1DEA6F2A081C2184E6DCE94A5BAC95D51AECF492018FE21F2DC7471FE58C96179D51684656B4A3AACD2DAA6C295381BF493AE848C21573A6F710BCF99C33C70D2542E7DC980E4C37DFDD6BC1C37E41C14F9966563300C17F7009A7AB344CA070752A24BAE942D70AC826038389A7BE4A37DDBB73BA2E5CE2A85F9699F2651EB8FAC9EBE9987810B682450A1F94A6A2AF5C545C74509F3AA824F5842CA2F18E94514800393FA391C4535B8C8A55D8D7519AC81C5A80973585E31E0202B7BE5144B67DD8D9973EBBA3CFF3E8B4EF14C529F0335C76E654EA33AE97C63F15EF3C32FAABE89E36E462B1ABD8C3FB645F94F1B3E6EEFE6CF34946A1811AD5FDE7E75341F52D2B6D61B5E33233664EB8F017693621CB2A0D0B6E6938F3E69E44CF9E829CA6BBA0A3E8EB130E9502E2345AB83D7AFD304C070FA126E44D7A8E98E6C2BB71306259235E57E26E4A581C2A3E6D94A3AB0E5125A06CD2B9F5F1FC0E0724F1355F4BBF7A2199628972E7280D609D0952B656375507FA53FC247216B61C893E3B191BB720F2F2713ACC4F977015EA082ADB3CC13F26EAB31BEA8BC7021347658A68ACB1A0B498C8F8FA8EEB65705676959746A3ACDC3C4EACA4E1E52F90F549B81F85AACE52408681E18A14C7352439E889F9DAFDA5FCE31BA1B6B3F3A36EE108765BB8DF496EEDA44196F9B7CEC9EF5A2DE092A94D2DD3AD265559A4DC7D5449A809C2945A443BE40F1B4CE373115B61918328CB8AEF08D6A3646CE45926FE97ABE4465F80ED1753074DD49D5C9AC8131965AB228ED7EEF703028F3A92CCA714A0BA39FE374FA9844E1DA950271328DD4FCECD4DA21D4F0D84F1F68DDAB2A38355EB54052BBE72565B18A716A790670548D3D00C9EFA1113DBC19E582820F93F536532FE57BDD1F04D56FDBA8B07401AFFF347DF41236509EEAB938F10A35BB2C13C8C93B00F9ADC8D30928FA4D772DC3AF073570E4C767D1694616386E92B48B18EB62AE3D6196BF5160103C50A033E851A583D6B1F26152DAAEAF1ACE048B6084842A802E5CFDD7639ABB4DFADFC1153A67A895779239C22A948174245BE2DEA40030F51A43D705E05D7856DFB7466FBAEB058C7189154B8D3CB5AF438F585C990B22B3F3F7C91BBB438C1CF41E66188F8AD8F5BCC02C486158DD9B6689B1327E36B93D659B7F21D7291464F9093B46459E180285FDA4956CB79773E067C8696F975BD9248221424F784314DE8B7890BD20F6B12C0764C5C0EF4E183D792028639E9DCD2E18F280208616AF75AFAEE46A9AFA33C00779F774D88E41AE70F69C239D8B2297B3F18EF3D49080F9FF0A24B5FF2E24FB018E5D2FAD4556C762DCE73F9CD78BDEBE1D4BFCE89D0B85E25C2C30FB4725D7C46FCA86755D2602455293E6FDF5B8E0BABC7B9EFFE35455C570E829405BEC6F1B07807F351B4B97C020B39715FBB1D018A6296AFFCB0C5F59D17F409F25143AAB82EC5CD7B82776006D34FF0E87E9187B64FC7F3DF1B5D461F100F33194A971487B25C40CBBBB1E0DA241BF7F031E5C8D7E858680518DA65C61E7FD994B5BEF3EC70724ADB727B58693A18F3E9E324C9DFFE793BD97A0B459298FFA63D40562708F3B3F396ABF0C989FCD63A61A87472026E24783FFB7D9F5D911203B595299A34D9D46149459317492C4CC436BB6794CC90977CE837F789A34FEE00FE2EAE25F2151A7B5F9C76F779F87410D6AE7A41B26BDB2CDD7873CCBFD243033E30A12641ADEC75B0DB751241A5081E4E5C8F10C3BE8BBA2FDCF0E50DC51416F3F07396D385681A93FC041E9D5C2D9F8AA9BBB95B63A0CACDDD1EC785A3EB4767AC093C594DD450C706227FD73472B36356EA0B19E670261FA1AE157F0A0CFAA8275A14FBABE7A10F698F035F00E23DB6CA54283AEADF68B6565A769DB443C6F34F1983F1BECF26B48ADEA96885A142EB9BF69CE2DBAF66EC7F142849CACF70A4B5A1D9A2590B5782435F00B0586CF9A96CA234E6692FDDCF8ABB04693B22430A394466A48FE6D9DCE8D261A556AF96337F799A1A928012AFDA325832CDFCE4347D36704EC186A572F77ABA6B7850015502FD13285BBE08B0D69FCD6B07F379AD9AAB35081CFAA8A6B1666D017019F534FB5EEEAF6B3D1CF4F029E4EF321A3C47B0267B33B54F15AFEBFC0F1FE79C75B58D0EBC384B5A0E216A2AC6BFACDF990AB2DF45C94575E285C6626E9FAC82E6A5734AAEDFA5534E087A997DFAB8813A711F1AB70EE076C7257EF2EE4EC576D688FD7477DE5F9CC3BCAEE55EEE9E1D1CCA73A2B87E253D7E1AE90B9A564B890EB913880C971A9B49308C5239121CEC2953B1919CB6473AA59C56994ECAD2554F15AF5195C0E22D1D721ADAB8110EABB8D3DF3AEBC5F1E73029567E3F769787B0928DF17658A193A06679B89FB33C3A78834E7ED279C859FF7DC72B05BC2618434311BCD90BE90F23E7D193A8432E833FA2AEC23F2BAA4680BCF7B1D6794919CF31078847248DA1E1ADC03D257A300ADC5879210A8E065E85F170E67470F31946B2BDCDA525A9F1604B9610772D99409D3E74CEE6BF16EAC1BE852E70560501CDA994BA21C054F6C971016061C8A4D385EF5399368CFA7188B09A0C532A090DF87300951C581B1A90F52C0A21C962E5AFF670721B1BC5985B50465A2D58C93A50E22B91672F6687B7C7198BE04726D7D0FB1FBB26DB974FCA2E54C0E6B3CAE792EC69DFD6DA53DAA989B588BBBDF3FFDD1B436F34BF6CD669D564611107CC4D793CF74F6D27EC05FB5165B31FF14E3583BDC2366FE81295293B5B7F86F5B677DDBABA14AD2F16589283562EB176FCFD558DE71A28935091B44B7CDF309125BF5CC045EBF7DCB51396EAA1CF3D45E677992C630F62C3C42DB34FF9E63141C8BC2F3427C43AF748D9BC9DD56EF6BB26480F792229DEDC959AEFEE108FE2B907073A4C1C1130474A391DC6F68022F787817BF1547FF9F34553FABC85814A35097D33C586C839AA454D8FDA7C1A3EA10A0D233BA222A0CE3AA29353F8AC3BE05F8D60DF396E46D0224507DAA0D3929E74F33A70D24FF73BBC6C7BB41393A53273D2D78CB00B94CCCAFC82CE1A82AC724F3951D8613EB511B26CD17A0584AD52CFA224A5273775C388A12DDED328A515C832E23C33519697338563F643AC4403F7EF98135949A5D807E94744FF2DDBA8BEAA36FA8456C51A172437E19632A725E452B9C945803890C612257E1D9708A0BE011B24C0DC3C14036CBB9831529B5A981105B0DC62EE3D54948ED8706DE2707A82FD7B03C9553FB7F2A522FBAFE59243D30CD40815DD122621B1B31ABA7301A9CB479F273298266C675190D1A65008253CC8B26C6BED43122023CAA3E8047950F996E5FCD1010132B23C70EA0E0AA8C058EE009DBC1D00234F15F2D5E04A74DB7CD0F80AC2115D5D7940495BDE61B17466555F158B436D98787A12660F5FE1EAFCC1C26004C229627D4E75859C0F6705FD2A11D5C3670453654D7F0CAAEA1CF121FF692C5EE1F1EB5D23E9CE672D5A1DD622D49285392830B5C07D559F02C18415734413EC361E83FD91DDBBF5F65063519080A1DFA336EFF27704DA0376182A7D0BEA0905101FDD8BB9E1D61D15B7D28F8565C0250BF5BEFF2B3210CF2794E56B10295DB88A7FA721534334F77564F967F93CB9E3E84F7C44DC0BD600106E040D36F0AC8B166D6B99980828B8268EF9BB4AF519958E9872478DA04E0807AC524F60E41B6365F0585B78981724AE621EE7CA92A366AF3F7593640446AE4E5F1336A77E6648EBF43FC44F8AD20B6CBE211843C94F352A9216B5D331564241ADC8616963BE135AB8D39F09788B3EEACCABA278BF94136AAF048AF692C4F25BA53784FB5AADB6CDC7D3A38DEAEA13B8AEEC386A79130BF02DE779B89132F3103153F230E64881627D814F5C13EE339E9F7D76336CABA23EB79656F3003AC01CDB7558408BEC7AA0914D3428CC20827E6A0D5135DBA0DCB498BB21B53F2B2F058EFC5A6798093F5DBED571BB2899880C1699E98D6680A585D4D507A19EAC850DB78925F4E40EFAF215392A1C95F113D1CCD38681059959C9BE80E10DC287864F0196D4A3276F5A8D641548A6142916B563EE1E9D88506BD501685B01B97231F9C09DB3E88D5B6C4C15AA50FE684B20309AC33A4DD2115D4901128861283B14201E754B5E61C6FBB06216E1399FCD873D86723AA245FF3A8BC81DD0077334071618BF2B56FAFE71827F17F4C18A9AADCC61D40C4A7E345437DF9C82988423A38DF31011855A8CF8DDCB033502A1D2FA2DEA303763230E41A0A37AE4E5B04B15E942373C3FD6EF1A87C77D1B45CF08229E45404946F79AEF7C0823233A0168A518920A928FF99C348E62437E3EDA5A9AB064101EE7D5541E2528104BB3EB22DA34ED9EBEE42F80F0792064546AC727D460139CEBBA128C7F20B7BA1BBA4E2757AEBAA07531A02FF18045782ED27BCCFC00E5E334D82B134CF764DEF93DA9C61F43FE292F6E06800394392FDFE95EAC3ACE71B1BFE3207438D62B01791E25FDF82A3BB8628EC542CAB4A613A7488E28DAEAC292899BEC6CB5B9E0D1240855900B526ED458E221014668E74CAE2650291F75A0E3D8C0A672E9CA9B7F5A5C480F6C07966DC6CA88112F6212320C2B7B1581EE3E262026BF175DB2E609D57E394528034C0FCE05AAC07C3563BC3030777DAEDFD15E116AF3A60EC29623771945B8755C5257B61967DEF3D7E818137932E1D3CA3D0C19CCED343BD4ED74AF18E73623FE98DE4FDD69241FE012714F18DEEDB217B2EB66FFFC788962C3331DEC036CDC1ECEB64C319E1761412942A41F10E2DC418651312738677F153830B1CC1E375DED4B15B6A815101CAC7846E7039F9738DD95DB97114FD587537AE86E5EEACF084F0C0901F90DEEB8ACD4BD7701487B9807717F4595725C8A00BB492C35DE5A43945F4D90DDB4440C42137F781890B5F518C7C4FF4C43AD0DB69B8FBDCA3309A639BD364D36A8A342D1AC38B4D4912C080A253C7986AFA48A83C6531827318CC8148755763D03C0DE1106F1C81AF03176C374B399CCDBB26A56744702978AC99725B64F1A7F95B010CBD32498F18D656226954A60440A981F84F15834E7C243B2F902113664B8EAA270178AF3BD83155B3C605661F93A27DCEF84158C27B8747774DF077CCADAA6E4455BDAC1ACDAB7D538B5635CE62B9B1C58F7CC5B6A1B0DFF3A0924DE9C5B9AC0399CE726D4A6D1E68F412D3CD09FA8D2C550ECF0F240EDFD607A76B501114781B19F1CA45BC2C31E5F3401570C9E7B177151DF8D4563A4D4D49938637B518AE8B651FE4CA4F92D903C7774EA173C8E60CB4F38856463E26D006B6492AF9C1EADB9FD58DCC042DC92AE9C017E9C3E4EC7A0AABFC0C93F502608D525667E7486424F124F81DBB9FD527782762B5CBA2F601AE6ADA34213AE5E6D641DFE20AA78611ADE284FECF020906CDB188A88BA36BCA472DC7E7B818521493500B20AFBA5245C29ABB933DDD67ED160270A2C20956E10FE1A1FD363D3F77CE9DE39F67B29D86C0D6DB5E0EF0BB0C2CB26E20763A8E16A60FE5AF5011AD747DC207F635167130D7A85AF08A04567E32A54AB013101724AE6F23688EE3C4A1F51DA68E541B6741E7CAB468874649C066A837B377782EDFA9BF9BA7967CDBA4CC500AC93B9C7531AD708785B2AA1B190E49E71C19CD8D3062478311BEF7F6B6A2C273AD2342D34F7BCB53F9F903DA3DE3A7FB702B5DC1531F0B87F4D2EB682E7B7B24F8002D8117F1707E42C68ED7B7BFDAEA6F36C8C31699EA09BD132D4E1F859933FB566E3EB388422BB4F4D1A4B6AB0FB79B50FB98CD6EB81B16C456D9E605CEE55CA192F50C752F7F225823AD7A87DA17177F8BD10781784477D3DA7941B75415CDE3CEA6B5B4554D672867C0CCDAC783603F42B60D5E3C147AEE277183DCF63D7A300593CD2D0A811AFE13D4AF2E2F83BAB6FFB8ACBB2C15703665C3A1FEA1CBD69A6653599EC78E4B706F68BCEF81FB344324800A918411EB750E3E034FBF47F3CBAA59654EA84FB67D07A2D31057F537D983813DC2A858E8C7C54BB4887A0173E397542D7318A2CA89C27D131C9381036E11C712FBF4A1F706DDFD98BCE5CB01035E73245A8B6E883F5973A089AE864FED252C7D73DFDB2314645901CAED9459B914B8B19C046968DC82023A241F9251635D96A7CABBBB40C6D0A8853668740BB22904656BD232336A412C609C9F62923024F5E3E87881FEF4C6B36A484794989BD4D00C2FD93A393E777CD90595E61E9AC410621AD49C5BFD2F28309F8794B6E24A88735195848817A8FDE3726AB97860E968F036F252B2CB9164276BA64C2AAD2DC7FE58D054852C357CEBF33EC37629E405C21E78F46FF2FEB7E96EE75C6AC3C76C8B4DDA4400FC610DA82D7D926E3384E6267CDAB10FD87BD8E4B3F6ADE86FCB9FFE0366C0ED9D28029112DF9A0282BEC2710E543928512AC7C45E0620CE908F3506A35A8638E8D91BC4E57567F2A71FF61610172E7E68B3335D927ABEA7E8B414F5DE43D852340C9898FC4D94E628F521FE8CA765E068340E306D99BCD33B8800620C639C9BEAA686AA8DEB6C8B971EE3622DFBFCE80F7D251A7908FE2D6E62506A8090649C8461BFD017B332AEDEF430FAC415143D8DF6EB0C61EFC51939EA4D06F35489826CDBB41DE2CD3F28996C48D0AEF8B7E756D87F922F77C868C16D450C2D58A3A35B33D3F692E5CC1884FD10E419BC6E13719F352126E0B3D6AF37231BB2D6348E62C4A164F855248525DA95584FB5618B89D11EAE424670C32AEAB4681F4E48E1D0965C81B53AB12B5C9B5868729B2F1C2304AA28A48D2F763C622392FE7E777CA9F46B536E13E154DB114C7E89FCB7C5CDD62866D4D4B90BE6D87AF2A4FD72BFE8D003497AB69B9F91A7310A780D4227CC90563A6842E6E90A3F860BE2CF71C243DF7B429CFE71B454B3B1ED2DF940EC331D4E5621A77513C98B938A1E10825C4DD0758427313BB4794696326B57655B00837C7F08A3061CDA7CFE6D2949B2B57F1FCDE664BC97D6F6BE9D2B09EC3412458A51ACB75328FD71C6DDE71FDDF2702C15AC21887089DED54FBB0EA85BC8D3E4418079755A211B3827B44D8439ABC4149294D1F94DC6B0DDDE9ACB5EFD12266F8F4DF944A831C8B86AF9E4398386F35E3CA859C2918DA387CAA387013186A7A5ABFD36D444948DBEBF753DB3AA90943E35A7A45B8282D82AD4EC058443FC4B74B52798807EEA33186D1461CEC8609155E2BD1125B214315EFE0E8EA52D2CE6E4D6747A500259DEA2836BA2D57D6B5B87881292725900251599EE07BF7EB175CFB828BB95BF28429A2DEDD7951004F04196A4A036E970DB76E353C05B14F3D71471EA0C4DBEA06FA56B8AF580B469B5019D96CC8B83EBDC476642CCE776C4FCF4D5BA85B60908BB8B5E7F6F0340DB25E19189D03DEED82551C4DA20127F69A63EB15A822193AF845A80D9E8AD1C264108FBC2178C72A289FE687E712C5F742BA48784CDD6AE9BF31B26DDF7CE7B730BD361126A8B2EC05EF1BCF122FE2FF7F90E9CF2F278FE1652B807AD9A11F2A9FEF2F00F1109D05AFBC9EFDD838AC8D77D3C17BD24BDC43D4206020B63F8309A4389E7C31F5E7AC79192747CD52FE31BA852F95A2B9843EB6D5C2F45E0518AB58DCBF91429B83E5DE10B29D5549765885C76C481111D41D4FB37951A6AB9989D46C67B51842D8F1875B74069D791FB3F46CDA6DCBC9397C5A8ED4575CFBAA25517F23AE57893DE5C489392CE6083C5759ACA5AB9ACDC2C0470311C2C44E98C2DD997A13A33B7BB4C8818D1B3A7D1A06708A7B6B0D72F98A0D71F8BD669E348E5DF06BA531DD03A3352C18C7B1D7A9B0507ABC7E2896360247DD6C2812C4CA8F6FA0B9B634656882C129724A479F7B69B5C6A810BFBE5D5D41593F1A4EA072B39EC54297FBC62C69570B60B029C9D3D58F401827AA7525142144B7B31E4511A18F476D653AD28263A7DA17C089C61D6B285615F6CA7C689F781B67D7F99A7E1D7DA037148CF87FCCA8FC72C54AE6F82057B73A02CE302AFDD82D60906DF67ABFF6D6F75613B1A9CCC6B8AC509ECEBF3599F1012281A477E59D3E37FEBE55C7F3C2029FD695BA7295A17328CAB8C47AB0D6DDC0523729B3DB76036822332DC59772CC1725BA10E5E3AB4BC639296D91D7F9AD2B3B636BD3D6D106B9F766EBBFB0C2CFD6889439DCD28A79F7D7EDBB9F760B3435C140A1CFCA56C7B07DAC9C346AE128542D86FAB85BF534415CD20D24EF24B92F58BEAFA3E1D506831B21E170E3E666A7DFC45AAD04DA23414B70B1862CDA68A6252BD85C28318F1813E9CDB86D6872A207476785A10346E12C06C2D4414E5D7BF294C51B310C1763DC020FF36EA10A13A3A26B5271F18C254698DEAD54DCF7FD9C3ACE105768AB4607A6BB8BAAC5FAB479C088C60905EA212644266A1DD462BEAB44B04ECABB742A8E04DE3E9790A7070BB434587A28220802CA6BBB7502F0D90F8B09DBD676CD19DF9A2398186B423B869CBF2D58CA152CB0998D3CD8F34297B402270C1B5A33503E038162B7D55B7F6970D3E0FB18F1D6FE8DE479DE57359F501C6F9E4CFBD2C83D5BFA1131DA19E0230ED7FFB42E8D3B2DE0813576BAE13724FD464351CDC04530089CD5F73EB360CD0056DEB36BF1BD134981373727BB49C28CA977BB9A4FF4BB7166EFF1F63561DCC7ED341C104736C050ADAF4B1F327331076D313C3E5D08FB0FCEA5E008058DA12CFDC3C50E4F046E4585B9AD394A53C3486B0C994209A7560BCDC65469CCF36C16B9D8BD8340DE40BFEF99C3593816F553519EFD03EEBF2C3455727473F8F09D5829858D6487070815097CECBEE48F76AD2F42AB316C4AF59E6F7FFAB67A954DD060C539277B0C9248CAD6021FD198A3278A981048220A05F63E9C8E35B388B953D7D6629EA3ED892A83A000970FC703B51BA4E3624E4D72CB8A261BC1A4060E9C8D02EBC1E1EA2E5CFC8FC2F174FD5E2EE06BEFFE6D1F972697E9C1C5EB98529D09E7F20861E469B850B0844A535B4FEEE052959E499EB7683B4520D9368C69227DC8FA67222F6C9F83E6B26A70502E390AAABBF42C3E04409538A62820879C2BF5047E4BF2E8C7B667E5EA32181AC2AAF73FD73F6DB06EAB594768E3F0A639494F5E309A7D10C69EC779E2E7DEB9A6017C31281490720FEB14CF852AFC490C796878EE03DF5E567EECCC05212BC92D6660C1EC087B3191E5A1815C7BC13F501C8E24FA1F2E7AD66FFF0AB5CFA626159DBC6D11DE7DE7279D71FB40501EE665483B4B6F04DF234B55A31864FA3C024012D3FDAEE12580E357CBF53423BF6E4C5C4BAACDFED7AA579E0E74EB9BFA0BEDC8E2CFD0F45594F5BBD46944BCF37DB132D1FE6057AE76B65C770ED025472EC49CC9D834BA821725EF4A6381F5B7BE10A39954FE9FFA524A713269A184B48B2427ECF696CA6DA3B77510EC8E997FC68444C411D51DE01164C223BEC300FAE584839173F8133C9396806130946B07E2287CD84351FD59CCCD3925C33DA7A94D80FFDF970609885560EE95395FD9E7E76822A26A98D0FF40CE26B24DF5FF64215F18B7CD3F5B0BDE9B12BA0E0E02933EB2FEF6F4A7369B2BB39909F048087390FF3320CB2E5F9EFF02FB49E450E8418187DA5F6A03AD3F214543FEDEE3DB792CB8AF96EE5C2EAC7D1735953B09E1405C245AA72276E75A729F33C6C7BE9AB07CDC329B8C75E131B1AEEB1BEC9E40A8C76F3BD6A6BF644EFF6A9FB6435A72A649948FFEE168425C729239BD732BA51E6773682057389326C846CE75BB4AEFE1C7F2B74AE98BE415F4D0B1EFCDBEEF2896EFE924CE030CCDCBA0E720D9FA1C319C7ED7EF4A08847B703F5FA1AA60AE2110138614202B9BD1FA7642C1A6B584EEB206B381D690BBB8CD0E355A35AAF8012636158E12992649F3B8EA26F1EDA7A8EEA00A6E331B5EBAD667A5677FF148B34FC184B078972DE2A88768DF006B7754BEDBDDFD9F63441BBFE631F5DD97C8D520D3721ACFB67C7D253FD8F177AB95592D9453655BF925148E1F303E1EA11092CF6010C55E8CD9ABC83E03D8A10BB83FC156AA4DDFE9209B9956F97FD88873ED34B22533E4C568EEC9D1B30BF998608D89E0DB84218B018C92F3EF9AED88675F7D32BCD996575705F855538CB5477D60DAF86FC86FA3410DF137B8E40407C75D49CE0C45BE242394A7924628E795D0C641796965C60052386C97D6E1EFBCF9D0296BC062466127A2C2AC75E5E6F05EE419631EE4E179431B5EAFE6027E4DAD468CC739CB14DEB2BE7592E54699B84DF2CC8CE1C79D889ADBC3DE890F8F8F94911BAD56E827C824B2D5B41F57F6B8EA532DB2C257AF06662EB3EE9920ACF48140D61E5766B4D57B0B31DA88F43DC101A601A9C59B67D97582A50A0815573D213CF4D9AB6C375B8636F5F28DBAA6F4883EB8C8A6E92F1543FCE9ACA6E65EDBB2E2A2E2CA13F734B38ECC29DD4ECF12FDE2EA56218B4CF3DCC0EDA425BB451730A6DD313EE35C84EC8797058B797678F28C44E7422F2E222A0FAAB5A03501B53005BE78981C77FE606CB842C7D35238D6F1FF2C3C8BEB407C18D461F6E5C863A1B5213469F0FAA557C280473C948E996F6EB375F5428C26190CB062A39EAACC338A3D64A5658D6E8639E84BB1FE356E3F69A356635CBC140106A80DC2BE1949B4A4C6958A7F61E08D156EB8B9165E0C92E9CDAAC5218CCFBE87DCF7F4B41AFAC31F7D38C09EFD4DE6FA96DDAF70D56E26C3307F55314843E1FCD44D5F701E2CB5BB1F601FEABFF7C721A663D4080CA84B19EE601A6D2EB3C9A1ECBDE1B6C292A656F3258E6CED39599922E664EC940CE7C515C929DCEA3E486296FFB859282954AE81CC5BDCE50DFACC7334D06B8DDB5095358BA74EAE416D4EEDCDF6699B3DF268DE93170F36787A219F64CB3B510FEE696CF41CD65F37C2C9CD8DF44841D33A870D3E666608BB3E5E9EF0B5315E43191E6188D91722CF14340241E63367F11865C2FC9CD20DA0D14A895291D968DA9FDBF10D34EA9C65AE3EA908DD155B0C9C0FD03E3C22AA7EE85A23871A9F10AC24F02C1790C37879E4B1191F4409FDF02C96E41B302594950F841D7BADEDE515342EA981439F5BD1DD1E0B2E84F991B209B39BE740FFA4491FBDB94BA87F3EAE6B386D0B31519E49CA3077CE47C2E91FA123A964AFF5CC0C62A928D54B6875E67BABDFA8489EF0185C7134134C0AA1537D189BF127A18D8223DA07FB2994ACA1156BAC52FFF223AFDAF4DB00970CE5729571846D7FE929A73115D13E44AB84735281178DC2CB5BED1FFB778C023C21161FBEC511D8251CB8A919B9C8AA07C0D0FF05AB263107817AE4677341F9F0C39B71E7056147F754A10466E8AD797E9FFE63C9DEB1521E89A653FA08C9E0D4B91C4252595D145015F36C73F2E9557C399D0D98DF8E3021BBCF2B4B443BA34DC68F68396F7AF93DD9243360834BD093EF51500871E79611A0C55C6A04F063B377E38951F9023277409A2CF2B488C3DEEAD6C1F1C4B2E769206076B5E71523B9FD0D1A7595E2A4EBEEDA6EA82A6B18896BA0F69DC806092A9071BBBEFDE515014FEE1C1DBFBED5CE147C06701C669841EEC52D3A1580FC71242E646B5472CF62EE34AA45950D5EAD26625804FD064C16FF1784644B6CC3304AD09496ED8852B842D550E998141CDDB076838423A1DADCD8FBF6DE0F23D1009DC01B5E7F9FFD6422EEB053F10F4459025BA3C41D7EFFB59C88F9EB3133E4D173F0C7371F122A2C14DBD78EC3D60498FDE8D1C1BF27AE6CF483C56B42270477D3C830CE8148322A99079986360123AB4F23D7F0C7928F16C37F64648E27E308783CE748335D201AA4D70BBC52B4A4CD5CB8259FF9ED6916FEFC0DD369B71F8A6CE855F74CDE7AF9D82DA5E6598D12F2698EC57737C27EABE3E8BE2597327FCE23E6748259DB16C17F8F5DEA1BF90A3217623E1E17DA49AD96D96B45C7B43DD85E88A73515D11860F7EBAC6BB925E139CBDB958307F55E15D076E21B2ABA2B0ED265E963A59325CE2107C2244B329B6F7A216F04ADD47A5A51ED036FDB53E6555D49C286FD216A54A9BA2D3D249AF2BA1E3579579FB008BE809BCC13147D0DBD99B3F4B9816FAD3084D9361CEC15F3518C5D93750946B79E9E5E63EBCC1A655FB13B1D20858816E585EA8DC469595EE057CFD8FF21384F6E53C577A714AE7E55A67BECBF0F5786C041586167170EA3E06F3A8D94B18094332F913D9F5EBE1C682615C4D994FE5A6EE606943DD547EEEC7DA22630302751C8597AD6743B9939AF2F2293FBF11FC88FB8EB741AD11214E2C9593463FA3B4C50B64557F4D6D94151D1C3FF2D5EEB4F817F6E52E0D194FFC4E18EA11587B90DC4DDCA2B78275A908C4FBC880893C278EAEB5FB4713744CD563BBDC9361A883AAA8FAEE50CF40FE27F83BB61C545A1E828796AFE1512A6893D043E809B451A3455334C0288489D0070DE737F8CDD51748E71A67842F8E6C3F829BFB758F43B8697E1E4EEC71303C1A2B5EF8CC8CBA0B22C91336528EA6D4372C9729776197033769D9DAE3DC4318853F2C6C19644520EE56F83AB0AF4204F17F2D4C73FD60A87FB9CFAD9842A18BD30EE3ACFF51C02FBE55E278AB34DEFA65A2267FE5CAA9E0AA4882A12D0E87379F6EBB896C943F892E4505988DB7E9DC2487C97E6B15518C9423088E3B1E438E69195D286A744C7EEE97BBAD354CCA3B92980CEF58AC151DF4352BCC4D4957F164C2078454F22BD298520CF3A48F3AE2A361C13D3E3288C553A50972E55682C0728CF316A71CA1EE71B64AD18EBB986A9C212E89CC77874451593F81D27589AABC8ECEF675CD45C681E9C7AC9AE7BFECDAFC7496BECB33E7E40DA402A3112732E350C3F358F49C04D51F6FEE41826BAC10F7D28A998F05EB7A9A3991C9D31BB89F655323F0FEC2696F59BAF886C5A740FF58417BB9144448503008B753E5DF120B1409165364DA2762CA430F14D56F952FBB1486D22238C581C397688F830AC7DFA13A2CB859E159E356446F1CEC638090037C9A8DBDC25657EE7EC2CDFB79AF7C62F5F2AD176FD4BDD7B555CD31E94E5F24964ACE98F042888DD25A3C0A7DB1AEFB80AD38234CD29C580A71E3C5ED981A560C433C5539F13C7A2D2A11C0DB3188BECF512293EB8C392470FED939A5BD6FA548743C9CA9A617EA8B1CE9A15A8E4FD62CC2B690C28A3DFF6765E20D1EC036883436911D88920239327E42C3F368F9057C2DC2BCAD3FBCB5645987CC3C448D7FE1605DDCF15246123FD32676F339D0C3C18F7C5F78249F15D3830E538D75EBB82B6D3A6A4BF114D4BBBFAD6E9E7A252D6BDF3064D9BAD88E5BDD2BCE5E342BA049C481DAA001F562C2563EBEA633EA89882437F6EB57B7D6671A4913F971C00766FAC0A7188F12B7E4537BB5728F5DB9528467FB51BDFD96871636E9F3ECAC5FBEDA6559D6CE350D42373DE743C479FB6C7439C0EDFFEE96E5E3ECD8EA5498B9463AC3C1E2411672306040F6E396A122F11BBEEBD0B2041F9AF3093612C8198CB9569FB01F2D83D2BA0877098F7DFD88A22111E4797A8430414DB84280DCF2BC78CBCBCD284579B32E81970427EAB1579A68DE5D9007D5B4BFEFED5B399A95C9F79ADED00C17ED1EA4E14AEE6D19B0E06038046C75F6EC19943095CABCD38914B37D3A1D6F176B82A0D1C69B9BAE26B7567E8532433AA9A90063CE90A240D795965FC82853A586FADFAD4F09A253613BA27A13346A9EB3FB799CC7B650FC0EC3EABAAD8A9CBCE843287C234F32171B2DF9D26D7EC34E10E7FEDFEFCE0A8EEBC7E670E796D6019296314A79CEBA4E75953372C83A12DB5724CD990FD7987FB2FF6BE248FFD807541317650533CC39D0181F7922B2DB4143EB3BDDC672D16CE72320CE2F1F5CF85EEEA51474A7946746507745C5FEED8E41EC7BFB48FCB2C9E0159980BDEAB0102CAE11F9FCF62133B916D717805B55C2F3D3987905EF8EE84986A235CC27A97607B47627DEBF9A0D7E0D36A5F6E14680ADE71A2348ADD159C04B75BEA0558619EFFDC39F0F5726F28BE105AD5BC6DD961ED6157BF23EDC8427BCB40AF48091FAC110DDFC13FFE371D2E648D81BF85A6ED98427FE3357B5BA20080B8A345C38E2185EB56A861CA1C61927385297F1BA7ED788626A322606947AB7A954CA909358C349DCE56B9574065229C5EE45115B6E8A92E805B287DB71C2CAD0DC4538FF3E6040337FB890515DCDAE1AF8673C8F0EDBAED64502AE3C6163257E2B5B644409D0F701CF78D987E34C74EFB6E9D3DD630833936746072B46F1E25B5F4CB8BA0F6FA347C832D8DE7C6927B917322F55E662BDBEA4D68367B45415BD655EBCA4F8C70BD50BCA6BFF86F098CBACBEE440CAA5B421B67A0857FA0DBA013CC16F1A0B91F8993E7B9A90A5A75DC0F942D8B6BE38A48706FC399C928A11DAB51EDFCB4D6CDEB262847AA215A6167C535A5A3E7F9D8AECA4B0308835519D7FC0EBEAF9B297764971FC66B2854E87658EAA10C95C5863ACD5F70FC8FB2334A9FD08A34B2C598D8659B6064CB2F19915B66E1E725ADFAC15415F3C9C9F76E91D4FD968765D78CEEC6F639391BE4A4B27309195A3E4B50654C835BFBB665474534A82930D29DE86FF3E471A0761BDFE82F416E81526D242B3E69A68154A08D39E62F2FD0669F5170C767F2DD5A300C5BFE44FC515514D5103BE8248B5632D2C7F5B0345DD524CF3F0DD981014D343B73B044997B015C48DDBD168758242265351012B0357C639D171BABB3990D68762697AABFDA415E4D80C03F25069DE01442E39066CAC0096410BCC7B0D0B865F019E451D5131F839BA56859E878F302ACAE79E4B13FA4A87D5610AEDF3B7F6002A5FC703FC51C28B3F836E150F1202A16A7376C72E2A94C667B3F07109830875901C40C0DA6610E6AC713D2834EE72A8560EB41FCA1437028CFE392AF233FEFCE6D1D76897FF4F945D9F551DDC0686463BB67A2B823106E2A3210FF0953936921D3CD04DBEEA5C52A050D8F8CA46DE7DA8DEF33563160C949C8319A672D1B9B7BA551F87898D637A6B7880C92C32F09445D43E2502E87E6B0D711F62F42239620CE388517245A90CE09659A4A7159BB26378A9645289DD10640835F2168DADBD12AB1E1EC5B07B2F8662227D294F382AEA428777AD141DEDE357BA5DF5EC958AFAC533C6B5F21242D570A10B049626E50D330B23D7E1A5884CF6FA781CB37670C5FB7E1D0E0EB679D008602030970D018888C58539B2214B50608F93EEEBA199A1C2FCCF8BC5310956BFA3F0D16E8BC64E0EC36707F09B57CD0237DA6B09B1D41BFB7185BE7A42A4A4294FB5525840FC43D2FEF6D1A09174E9BEE46E7EE2590400F7273A618EA8151005FB13C7AF55E50F9A1D4DC61B10E81AB997D05829571555DCC5A12F279031534C955D649C6C3B5B1D7BEAD1338C7E509AE50211C06035AE4DF16710030544B714266ADD502286F0EE057E0654F040C51D29A16FC38775C0D21EE0FCC24584D30667D895441D5B7B9F5B4A99408546042D46388AAA869A9DF4475AF05FDA81F6F2F7818D9D800DA9E63EB544D6149E9C8A032B27FA97428FABC138040E0D80B90FB4686BF4DC1DFA2D2A1AAFC777C3FDCCC7F906899E260CADD401096A9AA209425EC18058C9AE6522893A2205806881EDD38CEC79CDCB4274E46F8AE96484B0F22DA447F72B0A20C25EA17983E238F82D6FFD1090F337FFC96491CFD2931D211190B56F38EF2370FA0D057B440549810417414D88EE67B2D7FA6B2B49593E4CE4D1834EC1415EBBAAA15CF3F3187719C6272B7315585530517244AD24A2CD41A06DEEA21F2E3A21C83D7E4CC986E95EFA73DD259E9F857A60E3007169153667BF84457EB5BFB57F2AAA3B3D26D682BA5E29C7D30F950E59556F185106A9C758B47BFE54A184C8AFA025012877158E810D2D1238CC7B7C0942E3663814F0805EE96FBE3844BC239B7DBF70C7FD0EA9B0EF6B384BA3B321F73753474B50A7AA5D7B6ED3D0F2159A7981634A73ED2E3D1C057A18E9DADA0588C807EC2A79FA0DD5213150A68DC9FB710BFE0BE3D391DBE71052BF1715CA02668673C48FE248508777B6F4ABBA877F4065122ACE6B9840F01A2745C4E4C2C2C2533B4EF6B340A981B65D3812FF21410AD37EADA742F764E611AA6B332FFC79522E09110D687313342D6D784F03215C9367AD041E7F6CE54E63544CCDDB6E650E25BFFCF23C6CF7D74C186990A50764FF6DB7EA080B8801A2B222AB40AE73A7C4495D3237EBC1C59E40B0DF53EE1906DDA7046106262405BC81672C9066A07738EFA3E36EC4DE82392D95D7F86EDBFF38B46DDFEAA37A01B65ABA8A2390926BA46846A9779C25A25D50EBF8734FB8D82C07E4465F90BD7B5B2CF6D2D429D49120BFE897DD7BEDD286C591F91BC3CFC49B3E15AC417FBC3BF2ACB8B4AC361AA51308347F1C201AE29F0B01806D9005D12E8AED9060530AB7DD7BDD785A1B42878067DC60D06B928C8BD8AECAF152EB160F4682E53FC7250304072DD28F3713361CDB7ABF7C8B3EE40D09A9FF3EFF12EBF22A8E6B00A19D30F7B55CB5DEDEA43E08C401C045544B4F01016724A1FD6B3E5DC91F1F3FEED8F52515D38A70C8575D11942C2DE4BA58BF934C39D9C491FB4C851C87392A5C35120A6CB6E7B0C13BA0B90DDA94C050C862DCB71093123150232234F238CAAE0A9C5040DAED0437A225C885E752E365CF1286E6409C6CE60DB82484855220E8519DB6B3477EC190F0F22DCAF1193FA971B22A3A19DDB19D27030C197518FDE665DDA920881DE8246E6BEFD71ABD62F572836808C173270F2BE6F0028DFDA370AB1C5373945AC1CF45DB6C3D9D08F635030276C1913AC416EFC2FFE9726F5F0DEB98379CBD3E3040600DAB498B9659A036CB1BAEEF6FFBC7B0D5C49E7716CCABB1F770DF797A3906B6D223CD4646A36E95E44272F01F0F25136EA7E156874CDD1B015FB524E3250636A6668D6C99AA1D22F67F41E43731E8655A4CF2B868CA337250D0DBDB16EB5F49F6702314B0486E18EBF55BA55038AE067368306B070A28A991F4B8D22264D2B7A4F780804BB100E9F8273405E1A36133FDD8B50DF47418A43B8B65F81320DFF8A898663F9A977D2BAF8A66697DBF575D1B902BC004835EEA8DAFBB65A2B87E4D2465E57D7917A74903D4B9488E13821B8A51E648D9BDFF48CC73A51F6BD1E40B2D10ACCC6A08BDBDC63884C165D4AD71662EE877403AA98DB0ADE7C252A6726175606B8D56D2D116678752CB4612E0F39E05A8B23D62277B80C0B721F355DC34FD8540442D832E0483A6741CF8AEA5E76EF4DFE4179BC64A4AB90968F194F1EA4CA5F817BD2983AD3BF8B67A17DBC30FADF968B8F0585C69CAF60B449F7F026F5E6A662BE934F30077013F4D0A41F2BFE0FB5E32DDB3A01E00CBED39C3FDB5AC0C4B70EFFE90E67560CC977A2326CD1F4C6999123525F8358E8E5445B4D2B1D9B7C4F1FF1059728F451AB97C99B7AEF5C21BB750AA218B29A2F2D3FB85050396CC74081A29D6EBEF1C9558FDB9324CF71916DA9392E8390262F3C956ABC6EF963754DAEA19BF47923B5982BEC30886F7E6569F0030BE280710A0C5B63C6327DDE93BEC84EA9CA00B56270B601D53F489AA2E9B0D2F38DF492660EC4D17496B4E33DE6DF9FD80237266174EDEAF5561E68072F28493A59571003B71385C0CE3978CD9E033E1682670ADE697C68E125FCF74E5BA0AD21065D37EE94739D270AF205ACC2EFEE8A01E79C98D5C9FEC799585235F88CC0AC678656F44AAB665B02D926CCAA69B7464B7A2FE4AC379EB95257183894184A4C2F1E88E915C6706F124147431B1756788979F955DDEE492F0C8C3FBEB4C34E27C800E103C69C4ED3280DE0FCAF1C4D031BCD6768F0E4822E90F955BE853B78CE12C811012CF6FA17BB513CB34A4EFD1E3E3B2CE1403BAD99803399B161C338BC8D23FCC3AFB47C90BC83D23BFD012CD115AB6724524D259509113183CC2A7D5A6BD46008734EBF01237C236ACA99572B2437F78EFF239C0E19071D2EA03FD04B991698391556ADE6A8AB245E4E205DF3913E8CD2940CD0E2E1686DA10F79990DA1ADCCD1C353410E77D8D37642A2BCF3FB0146DFFA6FB3DF23150239C65DC0463091573D1D96DBBA4EB93B76529AA5'
		},
		SiggenCaseItem{
			tcid:      5
			deferred:  false
			sk:        '088A88C778FBC5E4B91C5AFFDC21EEF6A925413D0BD01BC37B43A27DD0A09150308082D86B3AE1C5D15DD578AFD3DAB537B27FD0218F5BC3A6CB94D6A96DDFE0'
			pk:        '308082D86B3AE1C5D15DD578AFD3DAB537B27FD0218F5BC3A6CB94D6A96DDFE0'
			message:   'CCA652DB6D5392FE48C2CF1C8868741A25231DBB7997A3511C6A40FA5B77A130ACE1D6CA88715C22C9282BA3AF080B3E639270799E6502A270DA4DCA755B2774657F2593A7D8AC969CBC217B39142C6935B55683EB06AFD1757EA23407F9DEEAA365B7DB7240F4BA155B804E377721120E54C45346CBDA1D5A97D49B92C1F21C0A58F25B273ABEF9099C4EC5230A69491A34F6F916E84296C0DE16303AFD566321A358A0C03B47044EDA3C88619BFB71C70E99E82513C063F9B3966E3F0CD34525B0601F7B3058B31C1B0DD74C3C49574C563D0D437B1382C3D4D119EE63205CB188C5ABF248C7041CDC6339968438CACC85D1606885CEEA5B5367433574907F54A45B840616DC1EB6A59311656FD62B18068D7EE375000C0DCCC1CE677EAAAFEEC8A86CAF51D15A04B5D56892DCB61D21CFC1DF247E48FD100AD5D870E0D48B0E25EE1B8CF8FADAE6B2FD2C721017E3A432AF3B0AB9D4DCE43564A92BB80D01E14879A9BF5B4FD10ACB99F95B2D3275B301907DE1B6D388CEAD76DCC904A67FAB585AA586CAE535B090F1DD41A38A5B122DAED237B85A3CED0074A5900062FCA9DA9CE58944A362D4C8363CF2C188425307DC2B00505A483DE3EA292CB9FDE7CCE39FC9E5DD62EE59AF239201981FD829A05F8DE72FE049A482C2EC33FC11F75A38D41199B2E3B294C45AE199FFCB00D01E263EB1581FA1F5397CC990F7B3B390BD91CC98EFF64FDF10E606D0D582204B52E4E6AFA1B4EC056D019002C2C37BCB2AB71C201653B405D5DF6645240EF7CA7E8B53727EDD47D9B1E3ECA4FC25BE772B2BDECD4D9FD7A656648CE88E9EE859A68C27813AA6F6088469BFEDFA0B6A62C8F4E30D679E57A60C8D1975E5CC4370D1E6AF6688876B0E39466BA445E43370D972B4D20FBA4056F3B008A5B5304EF00E04D22E7B44D57DC6F2C8A8F44A561533CEA534BC5175A3152BAA5D04320102EE5FEE9BF9673E7FA67123845E55819E0E0CD8B7323D50FD9FCB95BAC37CEEEA7626FE75E864210C85D8710C4E146EAAE56EDAF21D7828EDD5D7FF1A73C457187E7299CD00670CE8FEF52F5B2A25D49FE5097F1B956C5D10F3FEDCF54C2001B5339C3223B454B3658A6F5F7A881CECB1CD4C3A757A8BB5B0964D22B3CC96575D70B87817D7A2EB207EF9A64A1DF35D15B2A98CA37E716EABB30AC5A075325E31B97C6DE6329F5B59F0B8E7E83769BA5BEE97E62BC711DADD9FAAB632FBDCD965E1DEB4D84E4BAD98D454B4584F0D566A3CC17C4F97400F6D55BC32E0382FADA51136F58DD3F71C6AE67D6BD77E309AD18AEE62A981EB9CD76B87D06BB694163F2B3388E9DEE1599F6AFD3A33187AF52527E9744E6FD9D89A20D46E2D96876821B183527455C2BAFF3DD1835A85BCACDAB567F21FB6C8C37DA8DEAB99E09670ED57C0F0C455AA8D1A082A1632578179CC6E4FC30775C0E2A247A71FE2DCC32A5303DADBFF881A2A786E68DF986A0B24C7C1885D0AEA73C733BF79DF7F23FB83E8C2813D7B493A54CB5AAD7B3DF3A11B272642DE60ABECD540562439DDE68426E9A5D33A85324B0AA0E808F7BFB41D58F956C60349E528BBFD076FC754DB3DD4526D305A4C9B72ED2A8BC48866EADCB01D79151BBBD6931A001FD5F81F769665716FE19B653BD10E7281DADCFF28DBD3FF8F3EEA40AE43340995961DAAE46E0568C4B142BDDB405B6355CAFE0B9CAF963D80DD8E7BFF2922B19F77A59735643C80E579AFBF1853DC1EB9E96AD1F5D3803B2D520F20EEEAE174705A10B85E154DBF9BF4DE1DEBC4908FFE7D66E19D930CAF3004AC8224D774C4969A83A8E3DA9B1FCB08640283B140DAD533F863AE780EF403F493FA3518C700F661CE2B9E65C3F6E11559AC8710A4C4FEE19AECD86B2565C6220EA6D17C3524B4EC1227753FBC7020D1CFD4DDD517119A65776A3D7CED0989446A5BD5E3C8B0E937829F223E2A764CD869C574AFA9317DE38A9A2C1F5B378B3466A0B5084889974384870694F52400A48999B3783DEFE420631D6C5FF36EBE893317632A1AD5711C3EB29E8E51E101F6F9208D1AC0BF4CC9CACFDEB9A6D5F622155876F71BFAC416B374388AB8AFEF42D71235E991D3E1AA0E7E24DFEC2491773C573D4123D8092F0A1EEDA16A5B47EEAECBDE374D337A52999ACF2429CF35A016A2E6009E9E0DB54A821C0B257B44DEA34DAE21C5A7192258DBDF308E53B1272A131DAE3AEB3C5DECA3DE6655D32D79CA5E77DBF75FB3335120EBDAFBF95928E972DF53F40F3D1A29A68079DA6A4344B6DB2AE87C9B9A096712BD780566036D1CB9D19917E455F547F47691681B450E98F140FF6776E2BB0CF6374904840F9F37E8942079DB36F7DB925E5E56A6009F5BC2FC15063B56B1DA4B754EDB3087A553CD3868BAA1D19507473ABD27BC06814513798C2A626D70514EC24B713D3E164F861B5D2845B2D54F277773ACA7FF9C97E68B1946D72C6E2A60AD6C7721BD7EBAE76527599E67D02CBF6456D098D1FEBA396C2EBBF8FDB5AD75FB8F15DF95B47E480B7DA5BAD604144712438CD9E326F0C34B0DD53BC6C6640BE12FA27C173F03F130B4BEC1C10646426A82BF61C08EA49D0C2D1E98A5AEFDCA3F67C01C467FC9D1A44D6888C4FCF069A67BEAC391A372A24CE8FBE111A73E983D83BEB270ECBD554650053231F086070F2F40E4473A4EFD19310904D40F22A97F99794B04FF99E75F32FEDFA18BD355ECD0F13351BE31B6CEC3B109D31D87442FA6BE054673D8006292A278F01CC0CB3ADD215B5451503E9EBFBEDC00FB7902AAEFFC61570E320E2C4584A2FDD0758D9FB2054D1F32332B08161378810445E734A04966AA607D402A408E877D5854B23740E146E3AEA2F455A6C2D44E5D4EBACD02FA5282ADCD80F8E8FCC12689D1CAEA62D6D0BE13E92FF2CB1377E175282701B4104F223F140E109F59CCDE94BF691EA34A7785506FDE511C9196BBDE2051B5DA55E6F2F06D35D95B202DF13A4B8362CF5602C6DE02579A033F9075ED6A31CD4A072918213974A5115587A809E191AD0684260FED9BBC046E072B6413462EE3C937D2CBF98AE6F566F0629A06C6A22FA4A4BB1C4DFA041CD322A3082FDA9573F08E6EAC113551C2A0730AF2B8902711105B3FA9BA1F7137E4E3014A4D876970E21A2B2ED7B28AE34D753BBE31E900D46DF08F984A788D1BBC455F9B199F38DC323BDBB86595029FF38A22483A2E7D447F1AE986649BACBED390C3D9527E6E70BD76EDAF2D80EF5776F334F73661AC801FB21A870FF6531FEB083954EC7893288158A9E7AE9CF69AA2F87CB8BB97C70CE5AF52E5A7EFC8675E9C4B231A914FF3ABF08EFE6D912F7198C177D85DB1BC362C53E63B6C3F180F571679DE0E8E5C19D1DA6A78CEF360CCEBBE25BFFF207DD77B5AB276AB21CD15685CF1CD5E1B30BD8176F8DB893791DFCA925D3955816B48E4D7FA3F4CDD90C9B5F3AF5FD22A5E48F77A416B6862AE7599FE543CEA830918BBC4F7BD632837C2E2613D37AC2BDE1ECF47BC5E99270DDC945E6784A0722AF32B5C8BB1482D90B4D8DA92763E42D30183F4AF15763474467540EAF4DC109D75D87C7A802C61137E5C33920D6E831C7F5244943DE70270A6DDB7125CACECE86BE801FA5BC2254517329718E7DA51FE889D97E0C47C8576D2D73DA671794615741A6D5F6C0BBA16330810C35ED547E383298BA2C26102D9476E0615D9594E28F6F5ED2EBED52713405942C755CCE5D8ED16FFC0A23C0B62492B34941FFA7076D0668F43AD34F983E92DDFCEC34C047B03250F49CF1E8F85399B63B75810401F2806135948E8FEFC5FCEDE31C245FDADE38CA56019997CE4C0D82BAC315951C75EA114C1F9E707A88529E24B024F5D65479511A9D89FC13CC80C4150908426421AE18020AA4442F4367EFFDAD544F00128BC30589C6CA9DEC1BF063BDB3D278504B890F350862277EDAD16827E83FBCE481D8DB8092AFBABD4D0A6CDBC2FA14C007E5DD113391FB6743A8297187EAF688CC36B7D8A27036289A42C6F3C96B270442E002DEB8791B49A18DF0D8C84500140E2646E9FE67A01AC4958A4EDBACE54470F1C6880F04BF0310B630428AFABE2491A2A0AEBF97F6096801E3677C3BFFE1D08BD3866991C6AED4F681F471181CA80D068ADB8EB5D054782019C5B38409A2AAA16AA7A2BB2B1C7E2F648FEC7E3981D7A6FB85DEAA933B33763194AE34DE39867E62AA99E44EF88C597621F103CAB9C4C80A91CD80111D5C049BE1B3B775F4515593B727FE49D238B905FFB7FF4FCF67F54C24392F9F1A259AA8E3B677B192593E1130C332AF10EC33C15CAA46A804F852696549DF22628656E9D71F3605FA15A0466FF43811D15A95F35B9215711F61B829CC71D742AF9E0568D50409B6EF9F53721B6609CD121EEB3C9C7EC077FF3BEDD0C615954D97CBAC69B14A20BC9732622C0A04ACFD328E4F61CF6F0E4C07C6B305B0A0E941BB6D86B8534C4B6170AAABAABAD84EA231AE71AF6750BB1E740FB60CABA15742DD2CF448B6EE9BB42DB6B27A8D824BBDC35EB707E3B67EAFB63D96FEF079183315292D06861200F8B66565D5F0615C1B0EA675B3D47C6C0A338A5AB7D75219938CB2DBD9AD5A6449129B845FB0A23A10E56E410A0CA4E5F102CA60FA5B13843AB526883A7241895FB07258CA6D7EC49484B5CB5B8CCEBA14ED4E1B26AA24CB7B55E1CE8536BEC6B0C9DDD8C6B9D33F2DF10B1F169EEA1C73BBCEE93902432D9949129D9C9CC59F93CC6A35994265D3D6871D79C7BE048DF38E5B5AD652931AFF671B2C8DA9C64B6AC2DD1B2CDD9ADF06954BCC1D4284A475A04752D8206270E7871334116C7912533ABC5C627A3E3AE1238B38C38AA2129B2C9906CC1986272F4F955B087BF281DE1F56CF552FD10EA7037C5E5781B08CE21BA013FE4721AA0A117C3388D53E5D81D2CA8407842E4B30974DEDB38'
			context:   'B67B7F53834B4E0842C140B48BBFAD28BE5629F5077AE5CA9731866B90D2B9863F985DE866950888121DA243B652C90A18328554F93C1F1364E5E88BD46125E504F60655C9C55B44AB2331268D49B080BD5BCDB6B7BE7D45ED26AEC1D9B3AC4444308C67D28665E5E83C1277820D3913A6C13F80A56915915ED9DC2FAB4380BD9AB434C75C5742FCDC721FCC4FDB1FCA565905597047F878F7E9BE1483425808096152A1D78F6DAB1BB0C89EE20D7B1DEE5F71034B8A1FED550C57C9035DACA41102D9CAF80D29C85D50E490344E844FB3C2722FE66A0AE32C4BAF0157CBFCFF40FCED675C2EDF608F586E566D4B39040DAF94005DECA1FE6936F9D76EB921'
			hashalg:   'none'
			signature: '99D44E950DBDDC7AA32C06D5EBCA496EA7FB75A8369F118DA9C26FD4DF37BCED3368EA7D09ABF73C9B06F715B9BD76C6489266E01DFD30C9749CDFFE3D8BA6FF7A2D0EE6FB49E696A393FA36DE6FEAB7F8D155571BBF751FF90E2C162C16DA67DDFBACFDFEE0A70CAD8152389E03A01875E13F3AE1268F22672A7B0C2495F04C2BDDE3E38AC2003646C7821CEE4B3FA61A3E89ABD1E80AE917B43C0C19EEBC9DBBF3300A8CF3E34E1F8308DE99CE15E8DCDAF38EB6210CA7A97389BFF4CA89C12FB872AAB6EFADD48DD2BA19000896B8BAF14A179C6502A2BBAAD7A81BB1EF408EFB72BD4FFECA20473DE12367F20CB05CA9C288DD44DE97104E6EF19A5CE9718CF2FF289A9639C5AFD5B130694FB545F3BA287E43BF429D079217722D311B28D917AAFBD46019D59F785E2F3B6EC5E7D371D184B9F27721829DA948D0868E0802F3B09C9148086E3D85B7D237FE826D40E56838FDA60F115EE68ECDD5AE4724CF1EB4214D4CF0C406665D6E073187D470D06E2F9AF385FF31EFF3A76F3DE5A8E154E24E60ABA581D7F8077CF3257C63ABA31C898DB8F8ED28A83313BD48ED0E8A85A5B70167CE911FBD7AE4D74AF6E159A689D60B0B588623319DE62F146A54810898642AD4C15DB3505BF34550CBF554A5D24C37CCC33F02F78F83BCB35C72841BF79B9B02947949A1EB86F1E4BA36E4AC6C8844A0712858511B55088709C831E79C194FE213009D6A4A090658B86421B65DE538589A21DBC539FBDBAFCD0AC8CE65D064D511EF3C205A44FBA7A42848E4230A6F598B620B8095DEBE9DC0A3208459FF90A4BA482F50A4BB5D8C075A74F47D8E87D8F69D1E99A84834827097525BF3E5F6DCF7A1B7E72E7AC48D886B3129603C17C27D97728B9838D6B9072E341303286F24C676017EE0B6A7B40F01604A45D68AAF4A3CB2CBC73179B78C004E0F096B45E937CAED2C4A4115DA0B11F9876829B1A87E2648017B666490919E77C4903777D72E57FA11D335054722961AB9B6D7BE4ACCAF33A3423AB9CE2E8CF8542BC64DE85A99B7309C3FEEB1BCBF2D7F10112A5029828F3CCAB685B1C4742C78CF2F91DD99E01FB88EFBAC57C52DFDF3D0FE3F9DEFFB1E2447689FCE1277CD5154C64CA972FCFCFB16E4D233B2285AC0DC938B08279F06F69B76420C4E3F24458A2DFA10DF6D9E9735487D38FF2330E942F573895380926F30563C66CF73A91ADC086E3BC20B97B0AFCC4625080A8205E9C46CA4720F1E2BD822C3DFDF585DB58B503536A021C7AD4868A9AE8FAC845FF6A4187EE9DDDCDD569DF11DD36548C5E01699180C1A5BE6D1D4CC0AA9629FAF5A01D433963E9F1B849F596564E9F09368EF97825E8BF88E993069AE68A3D751CE11F2D26E7D482E8B14929FC456265F5E6BDBBE120204A19D34E6C7E540FFAEEEED68AF9CBD479797A1E8F4D44BA67F4472F4CCBBE42F05F0E09CB5A55A15FCB5452CDEA1B60D2A62F6B20FC00433DA9B3CAB25D64791FF0B12DAA6F021F59C4EAC20771A595A596618D2862065A777C977435450782ECF67A8C5A1EAABA91CC47F7DAEA76B48224377F0F0A347EEB5C62CE9EF1C0AFA0BE8D6545808C3F7C410D9C6C6917570C17A9BC91DAB6E150421A9D3AA131CD9BBC2544988BBE9B2926F4465E1750667B0F8C75532A7339CD817A9A417FE742C2CCF727A085067D78B6CD663E74B85D287CE0C9197719D70F4CA80E43C45FDCCD2B57808B60AF3FB17ADD08437D4318574D5F5B068A59CA2A1A295F6ACEE2878A94775F7327B4A9703E1876651F5AF324E4074A3A0EEF7ADEA1606F122C606209F337E0D4BE618C1834E05AB33646B45B550D40CA743F3E68EECA4E709AFFF205B5764C17445D98DF2C05D8FAD2D82B7222E02235025DCDAB0A04AA8271AB8D6226708759E17A65239F796B29CE921A46B2BC75712BB497A8ECC32C6F548854768F33F1D21D769192833385B6724DDD55520461A78EB08689C94BADD1C91826841AD3EB95F892BAB81A1E8C9A1A4A23A455B3677E5687134EE1A6C6634B8E29B11C864C49B55811B7E168D6C052714A5E086FC26580B46F884A00751B0B96C76FF648033570DFF6236DC705AABC8C3FE4E5EBEF6165E3C109CEA03C15AAD7BF9C6D0EAEAE68861204D619D508EB5F2BCF1611EA9C0605A04BD123709D64AA2CDADF3FB93E5133D9B88E0EB025E67678F580FA20B33BB0CA80EC9574DC8D63810D1C6217B768AB2DE1E6116F716A10DA337F5BA315F34CCA220C5E5549E267FFB1B76FAA791065CEDE84BC156DB452196FA323FAFB937A2C00EB2BB1712DA8C5E867A19EF2353C603B2C1E45625E646305832F22824127290A619377A7CA6300654C67B375CD507AD8BE0373486EEDE3A58CF10F9A121C41C984BE9DEB7DF92313DF32078D8974A8C5ADAA58E04B74CABCF146E941E877028DE77467F564FE0F0A73C360A7214608B19F36A5A0E42DEF521A0A00719BB2E75ED2CA169F0E6B3F267C85C2F77195F488DE7D2AB7C7C2E690EEC876A440DB7C3E33355A814104D30A17A788D8634B79B8FF17A4DAE93391F7BBA4CE30975E3B5D2C8F21D7BF09F4536F9EE6B924F334BAD51D65C0BEAC6C767AE23C8D2FF769967EC68F0610F18D340A00EC40CAB353BCE2FEE96B0EC869869D1FB33C827C44E4E3846365C2D58F04B7758CC962D80CCCE72DAE3FFAEAB29C06BE8C7FF7F6532422E825B3F0E1368D9274806FAA4B02B0407CF32E684E3FC2FBEF6D1E1C0A04BBADDD383FA520F5DA31E03840843C0DE29009A2C4C685F5167DA16FCF3017F507E34A241E0ED0FB830977F0CC620676CC82221B33EDAF0D47FBB9D0A921CF76C22E2EEA332C9E30158C89CA8DD30B2FA7A67F33D16EAD7133365696C18F76BAE22C436749E63045F2493909245F13A87F1BA86881AAB3E68ABABF2CF595B0832AFBE70FB39E8ED960A3C1D7083544DF0A010307923727B7D311B388C699F4B60B4C09237C487C31EBA6CD199D6778E1FE7AD6B8E16628BA171CFC1428512015A9C988363E41A335F2FF9E53FB3972D8048EC5E3D4BFC9A6A13DC265C981052A62C6D95CC327817CF44A0D322EF52033D75294CDC9A63BA31986AFCDCF79EE8E42028F9F2957BB0406AE01143E64B1EE49162B375CD6AD87FE1EDE502086F61163BF5A75D1ACD719751D4A1115665F0F2155C77A6A51654B4055D3819AC76F325D4A49A92604CA8A58A136834617DA696ED38A542DC0FE7F6C8EA110AD958703449AEEB01A62F862247B2B8F026321676753ADC29250C9FED7471900F02C7D74E507D7407B7B949DD6BCA3B8DC4E29C7371768948A218A0FFCFD976811E6BD921E8C2199AC5BD5BFFFF0831367FF0C8058AAD0CCB226A7403A6F0FD36381CF8449767FE2E8C587D5369DB7F30AFA6D3EE3B0D15C3AE89E632BF4FDBD5D61A24933127B96026EE1DD548F442E476C658C53AFE5AF206EC8DD5D588D24C91FED0AD9C899CCF5802E34DF3353538F2EADBC5C2F49226A40D6713138D02B778F4027FD963F8F23B89A3A1B55EB1AE8D227780472BA59208632578CF7CA28253785FEBFCEFB80CA549F03D88FF101494F803E47A94F050CE42E3A066C94884CB5B1BF46735CBCE6390E0CC8A8C08D175CD30892D216C9B4836328BB358F0C9FC2AD936F73EC44D0EDFEDA47E7E202BBD9BBDA1945D80486476A9ED832E05AE74133C37B639C180E1560413BB6A434152C04DDBA47FEC31AD32F19A59B7FF5EE7D836E52ECBF073E69E6ED42AABC723A85D4CE822C7FB8EF38C573ED78B70E102708BFA51F7FD8A7D6FCE0AB4F0C702A2967B16331EF42200B5182F7B12257BAE4888E2354D11C2CBACCA2AB2255DAB158C788A1892AACAB3E6A6D698CC7351085095DE7A13508FA201177C1E6D7C4BDDC92AA2FBF555FF76A84329A9B4CCD002D7E0B1F5C237E3D975417EB5F06C00AA49AE6DF0B90B62AB789D7D9921250955DA0DD7DDB3DAA3E1D78209FF59097D50BB24EADF97CCE461171C6F7328168FAC4CBB8953FCD0198FA150C9A0E8E1DC52537F615233A8FFFA66451FE26A4B3604706CACAE3EF8B8226E3744D318C9D4CDE39E8D367D1FB6A68B1BA782E74E091457F2CAB390FBADBEFBAFA8E22AED36497630ED036F28F900D850D4D7DD97ABAD3F308DF56D6EA24F4C3DA7E82ABD5472689349313401479221D67E56104E9A0D0FB3CE90305393F2467B1DEFEBF96DC35AD4F15254D7D6BB1E97A1EB75DDE74429EFC2C05486164F7AEF2E315AF3326F75D6CF25363882C520C47DBCE310EC4658EC110BD49425443C49767DC8AC401656F4B395B7DE8629D7BAF611926EA291278AC3C5A94F1253599CDE2AAA6449AF195C7940C043F12F38DC6386180FA2936488EB4F2B74DB960BDAAED01C8BE1410B653BB3E90DD9D8927700AA053963C0DACD000193A0B6C6AC5AF024A352CEB90CD052F41AD1184CC68F73AF76115FAF9A46D4168C3EB53E7B2BF9F80B1C475608717E9146D7D03AA812DF38B060E723BBEF0B0C83FCA0A6C48757C9C87EF813862A2304EEC49A02221D908DEBBA5852E0B7705EBD5112CAED32BA0268506D6EA58349B4BF9A7FF19B7FD214FA0E0788F5FB81F195BABCA20806163A5DD2E688B3E4A55E942F3D63F64C7C4746AAD5969F44AB62F139E5AB3408F627D60A3B20182558037438766A0BD8FA45A78F3AE3D62290F6325069E8EB539D0196004B388E071CC62C411981E438CBC4626A175D022AD8447F0999CF3176A037357EC66C5FA0EA4B5B2CD1771455BAFA475AB03B4DF917DA3EB3C4756FDED89EFDA3A05EFB274E9C51BCB31BB9EA906AC8617CB05FE74B575D458F795A97B2483671C822DC1B8C5B53C52F8BAAFC6CEDE03870A598D77AC952B65500FAC671D2F10D362FB8484C976E3564E8098BF24938482F52BB58519046BB6962702483A182F17BA01BE444B245ACD4BF103707CA4942C9429B65591F043A0186BED3EF2A328BEAE6E4DC5CA9C31DC5488935871CCEBE66818E08531A94C7B8D6988203232518AB5E3C6C3164B6A3C9689F086F4EB10A4889F6CD6BD6D676123D388EA065BA46D7BB96F2564EF594A9FBCB96E4B0FE1F22D651629F5E60142EF7B4C0F5A9E93580709A4E3A4B21D0D5CDA2C8313B84201B42F8B89E9E4F98E840B574CED70B853513AD5D74A3C07D65196892CFB93ECBC08AF5199C74759E27A98A06D9072B763BFFCB2DEBF583F338C78BC26E8E0F3609452C431B259CCC4673D910F8924A9A02E9888582F5118C0D1342B5A2D40059F883D56969537E0BFB5A9ADE63F6AA1EC62F384C354505179028640DBD26888D7405E1288FD4CFDD576D47E624AFFC5BFEE338FFD91AC6311F72FDDD8149FBC8050CDD726CBEAA209AD47C7CCB3DC0BA5138D4D8DB1A6CAE6D22A1D6758C761CCC69412028F844CFBED7E6E502FD322AE8A35D2560FA6DEDB999D7615AB4C525B9FCEF9B407577406FDA26C7C2FE82B2A1D5ED44D9B12A5EE06B750C49EE51B67CC349A86C3AB336A281255105571D3BC58BBE8234E71AC43D475598E64F4BCF8C56FA408C9F06F040F599FDDC0D6C930044BB0DCA0D8C178264AA8AA4932264237594FDE1A50AA03352C563733E46C88B3EA13AD1B8D0C431F558EB8E6A7D7BC63367A8382DD2A540C0C24EAFD59B1A384343E5CDB10A397CD1B3B882213F8BCE4F4B20C576C6136F04BF7DAA0BAD3CACB7B8E3B324A62BCCAD5FD3EF65FE33414458048143EEF5DE72A2D9D788368FF5CF907BBF5804922F43C8BD5A6720C7261F5D44DE66F956CAA331642CA38A48D4C3C47C2931DAF927054119CC76E67F33A49DF6C7E03DB8CC55D3C5A9666E21208845CF5E7CF1173F2CAE3A0DED54A4D83443EFDEE6B8D2CB0CB3A161F789D484CC800C1A934E097D76AED41F0D9FE7D50F06FBAF2AD202D0446BA5C898F75ABEE926B4A982A945458A51A57C383C150A40ECFBC5E567A015F1670A61CCB9D4220CB88B7172FC9F7298F36E4FB2C39AE30530C2A795FBD8ECF1527B1BC04D063F399BDFD702292FA65FF0D05204A63D07046BF3B2F524FB12369227D258C3F71E9D1EC95734D8BC54E0945EC487F663B3D465C968C67CE1D04AA397E45FD58C9329AB2DC3ED351261B73116CDB86748077558CC716F1F7137B21EFA9BF198E5C86EA42CD6AE39FDDF7A83006941DEE50EB8455330DD748687E4510DF8D1B6AFBE548293A630B690DF040CE657DDD85ACE68F481521849D8335E24C7EE16687B4A3FE0B79B3E783DA13FC67F53435519294AE140A1C8C02B5804F1901835B4637DA75D4E3A7683786DD3F097BC514F9AD9647E009C4420A922106DC3742814ACA38D11F6CB10C8BBC4620DD3D2E84A3F506BB52CD846FC993440F576378F2B360E388C11E97985C0BAAE4A1AEE0371C5DCE541EB75864A7E9277BBCBE58897F7EEFCBBEF89F6B6BEED8123342D633C4DF7A4B13B43CD56ECB4CE07EBF8E32CA8722272BE8F7E69A08490DA3F3E1CA0FB3DF642A119092CFAAC6F785CDC69CCA02C2A5047123A9B1B221B0A6A07E1526826120E86BF07F536B279EFDADD31E2A3761709BEB8908FC9D751BF56495B60D88691685A0C9726A30D8A61243DB52F15F950D945D14128BA84A00B2ADEFCD72822E55CDE4AC736294003DF5C628D1BBD28A17A971D8ACE015958EB39435A7B44CC05E72BC1DEFA50910D8E6FCF8A96F5777D35B85B9CD81EF4670B40C22AC40F3686314F3826CF8B9DDB4777E8B721777ECAB84EE74FC8F126B6BD2812D7AF6B0C287CF5E0D6C64E2A89577A6C89BF3133882B1C59D8B9D6952494E00215966DDAA028F8B9BB8D38ADE73C5F4AA8EBFE9E07FB11A24FA372B8E132C6FF98389C9DED902562E8BCE16E71B993B6A565313BFEACAEA8D8C68454704831DE10D351FA659486F5E23B255C0FCB5DC02E6A535C64E50496E9F794F72FCB8677A9EB30A0B7A6BDC39B7E543200F1F5AA665BCE592649A925AF7B10CA71F4F5915CAA5D489B25DCEDA94D39096929F0957D995AE267B4EBAA22D0DB49961818F26C49C4BB780C13054F8EDE9760DFEC96781FA6DF28C2CF4CF11124C0BF148939038FA334A62F9B8321446DA7635B7FC20CD4943D1EC210251CC27D926351A7F3008E64E7B04D6309DFDA990B0732D8775CBDF6C61BB91F116FF22EF8D6C4FAA28AE767F96FA521B95B5CEB0E99F22FEC832AB1947834EDA3728B964E00FBA69F667FB48A53EDEA9BB31BCE2C2AC8F1D01294943CE4FBF7DD2B0E00CDE85A9434CAFC8A30C15087F8F24A388A3066816E8A61CF06E4BFFE18E16A0ED2E810DB7DAA2634B632544DCCB0D74287D55746338159C873F77610D8590647507C14B13A4B059FD2723C19D66C79239A8E307AB9024530D3FC4D37A8EB8BC506C528EADBE92736EFC9EC64A1A8A367BC9EA5DA752503E7E1ED9F6CC28E67C8F67413911EF4F0308F1567084B09973CAF39CF595D1EA48B008BEB7EF96E17DD7AACD15B1C37CFA848D39AA0D23DC75DC4FF7AE3AEEB4D7729CB23DC5685084FDF38CE8389FA1B2A7D964795A493E35BA65D38FE80D8C2BE63A6FBA2AD60B9CCA678F48DAE38B7404B73C438067C6B2852745971C1CAAF22C9B9D2B36FD5C9FD5BB9EC4FB3128C3A2C108EAECAC12CE4BC7F8AE1F16EEE5D5476909B3A2156E2C716B282FA4D0A0863310B2872EAF295F4DFECA03F72FD0DD3B57234D66C4702D6662384BBFA11D238AF1C86281ED65C288A5FC6F3071B867DAE3BE0D5B6428899814077F45BD62A9AEC2680A8494F52261E0722D914A96C86DF7D53C873BC45998BD67B301EECEFE91BE42C5951425E2FC0C6F942A41B575F3A28B1D6E3E0C8D3BEF66BCAC34CA9127B0BB0457B72AB54791926A845594904D29684F578084B5D65EFCC6755450CFBBB1D66CCB1CBECAC7F8E422F8D7DBE38985A0CC5105A9B4AC5829B8D1DC8C31635EC70C9420AA043887AA6F00CA5A801779E536F5387ED61F80D0C24CDD8C931CE79F75EA8A9F03AEDBF6B52E12F1412B68011CFA285D02EBFE6658331855C4F5FAD0B97AA56C46B0009EE113C484FCEDC71BF357126DB82CFFB2981EB045EE35C9E9A5A71AF6C68495B58A9F771A1FA470B8386EA5F8FA7EEA00792ACEFE733D5CB3B86B6C2EE506CB7CAA600CBAD74844960310715D68B6AD619B3B02F81927387CEC895FD4BE76CEA239EFC6999CBCD67D86A1BB2E3FA0EAC9629B0A54396BDF3CF247A1F1456F0E77D0238193D120EBF59F003887C65AE57E6379195799855A779E195D59E1DF0E5BE72EA3B7659AE526F928752EC0D63E84ED685DF21DEBD59555A087C54C4EAD002F74B839CBCC615C236D903AC72C537D19FC7DDB3A7B18DF50E2A9EA636066CB1264742974B7F4EBEAF71F443CEEEF38275E8B51082F1C3EE0B036C345BCFD405DFA5354099FCD651E12EDBAF1A647D5AB0880CD45E45DD9B8169A8CEC7982A1AE997442690F3C970A1DADE8DF7E916811612A00513C7CAE8873F3451E3A46EA80EADA1EB7041B394A52BE29BC919360D51A6905E62FB8E9CE8B85540D1F73E348A449225B78103FFE55BF8D1F83769E1BFD6A98214CAD86B9E3326F8C6D29BAAD594C9E81FB57FFCA59BF5A96DFDDB1E8591570A4782F176EF8D30EA5997048D5C0D0B405A64B4B21C6E9A5DB7957717636AEF5FAE38B5E10B0730FD9B45598DE2BC513440F90DB8C0F6EBBDF5730D9707F0A6982AF47E21A68DDDE7C5A279A08D826031E7C78829CAA924B5F6BC99532339E5B1208233AB48821B262EC0A220CDD5F39623F89EA5B627803FB2E201300F432DDF447B939DD0CE476791BA78F3ECD8338CFB03BBA364BD7D24FB6DE5D86D3CD19552D325D442A3BF365989B9B0F8D750BB9DDBC198FEF684D04BC6C745CFADA4593E789798817D70B5A62B4BA8AE6399664159F807713DF6BDFD51C2DE7487D5B584DEC5FD08425BF5B848CC1059702ED798E3C72DD485D0394F42ECAD299119DBEC9FDCBCB4BAF0B9AEFEEFC30938F79D7D92841A1627CB16ECD04E7CFDF46FE8A5B3F3D8331D3E72C96FFF445B8192F0B3BEBE1E0B1F6BE49129BBFF94293F64AC9AB6AEA864E52EDEFFB694DF82A1D60828F2837257E7531AD3DE47C21FC039125D24DC1C85DC7B10E10BE0155FB53368000D01F1ADE317FB779A6114EE4E65EA3EBE5C5D273C99CB969339AA5F439D862982898B9C3FD33757D8F0D8B9D1E7CB8481ECC5D3D725522D9515FB04E95F120CBC296E9DFCD88A400049B45145F9339C7002344A672E8A7D5FCE7FABBA0B210AAD5398090F31FD28F7692839FF061817BD455682369ED27779552F95A8276B73ABE258D7352FA8EA61BF9A3E94FD87DB0002DAB2DCBF4E1F47F56DA5559915F38028956003C49F36941FEB03BB79E9FE70D9D6B866E5376D6082CD28682836B7F04779D3C14B39F0667C92401C3FEFCF419008FE5C043BB95D370CD4897BFC371D93F54C45AB9DF92372FF7347D49B83D7F34A6521EF3631F7D285B91B958374071043DA49BEB7FD619591FA236C7C207CC094CE97EA4AF1F4A84D686260D80F8D2C9FD2DF282DBF7B48439D9294A16CE359D9692845D457B7FC9C30CF1C97FD6DDBFE888F8DA71C0306DF84D93E8C068BF6D02D9750FCB572A6F94B7B198A41677F3D08B1EDCE8C2E716D0AE0BF1DF07CCB7CD80B18005048DC00EA2A4857A632A2264BE17F4BE11007E963EE60F11AE7E8E5558D48B9CF804DAF2CBC31851D022EE9234AE617A3099894F120BD545F4899161EF2B88697264C34F4250A929C10888D3E50AA60686331FB3094B849263FF1925B9D84E257BC1CF955E8A47D568363FE9EE3E3DDF95FB4026513C9FF5CBC839077980FEA4A200003306BD95407D1F47105CCF51C59FFC0FE206251551753B0F7FD2AE46CC620C7F794A51556CC2D7E41DBEE35C0393245FB49D7FE6D90EF565C5F5CF771BD666DC803E34D9D480BAB7A80BBC470E81C9100F9FC932382E4C26943D840CDF4D60290A79B9D59E6696467000A5F71D2E543EFBA384D4D073A23244B0EA872CA5A929235C427854ECE330A5B66983EF3BCBDA042E265F9BCF10498C34FD6640F525DA685CB6AB8B917257E1EA27C00A63C2BB4D5F2E0B2B8022830A6C1BF0AEFB310AC0E4D6D9E0BE18C30A2F55CFC7860D099D1257974712A5046710A14E36AF8DB90365370AFFAAA4314321368E8EFFC46C2E3758171DCC1EFDBA3F633036A23B1078FEFA41EF04F0827C39F5FADC545AB34929115CF4A17391062A5F1647ED7CE77F8DF3D777BC6B44276E9B0008CD3658EE09E8A2DF76208BD1085BF3FF58222D629CA10349961EDB6515430361E7C8CE025486A4F0DE6264CE95A264CF502980DAD7834952374FB370538A4D11AD375E5FE3CECBD4FE0165B7180E4130A19B98342B63BB2E784AC460C57D267EA7811E1097497BBBB3CFC26DAE946B5CEF0456F0C3CD464F540D6771101B690A603D2A21F85438DEB685BC8963E395E0EC3993B2E18998E51F51BEDB551435FDEFDC1BB66B7755E2E49CA5AF6CA541A417E26BFCA4DF226ADA2ED2ADD431A0C05EBF35E3E8FB0A7F731A3D45BE9E0D763FE247D527703D89A33716C3B8D98FEF04B0876E96CF2C69DDA4513B945AC47F7635A72F6A443BE90582CB862C2AB746128BA867BB70ECE50EC97F1AF983C2C81A5DB2CC8EA3CEA2D21C23AF983DE2C02227D1947150DFFAD105430707E378BAD931CE372BA8B893C979E8E49289A939002C7DD2542B6897015CCB4FBF6E86F97378818BE5FD1682BCC3F0A34D9DA3B779B7A60C31E7925E6099EE05C872EAE123531F651DDB2E761F5AB55874CAD8225E5511C3B6704C97C1111CEE6F9CB7E6BD632C1B7ABAF811D1ABEF8D8A95B5478452D7F56750B4528B39B5EB545D34E7F402D782676407ECEF02EC2CD19774CA9EA12B3CF084B86C7BA3C0D58486A2042FD5F24F7A30B0F0F45746798A913DE5D913D7FFC43C08D931EEA5B272C8331B3CC9C8BFA42BFBD7D4AE2221AD81CFAA93549E1C58B4DF136CA515108A3F48F350322DF41DF87DFD199E4ED213E15B85B8831ACA6DD9C91CD3CE4BFADB2A29FEB92571C3732D1C64FEBC237DD53933B410516268A8239E89AA76124207DB1EB26F052C660276E51FE878379AA3C3A40EBBADF46DD7AD534FAABADB82BF84B0FE93D239338FB9357F093FAB72D123EA0D5950B6500DFB1F6208C60D4456C41705B51C995F3AACF57AABFB924C275406BF7252A0B85F8AA64B235E8A2CA6A547B62468B0D5489E418457780FAD6B3C45FA2EE03571796BDB5EDC9E7D6A3EAE3A91C110FCCE778AD203EA622699A6F1E20ACBEB0925E3635B200669E6D6EC8756113AB99546CBCCE256FE7028228EA42D0839F05F56672E1226FC819BF967223B40E6E6FB220026C717DF082CFFA51AA997A0A51452B5B9A03D9C3E8FF80168071084EED7FE15F15BDAE425F8810F39D4A0901CCA374E469127A5F50F162FC2657BC88EA8D77925544ECCB0ADC7A9BC370AA77FBF79B60264B3005FED46C1E5CBFD83B13C3BD536875A14544402D4C131E09DF4B5A9A7B18B98647591FD18D91BAC93F78C7A7A3BC78A6FF1350F0BC67FE2AE03F3419345387E9785E0AD12F1C7261EFC30C872AB247541DA6F1C3A4A5134D20D932227AC515B880B397C46E8C2CA7C731E5F4EF7BC035BB91ACEEEB97CCA103BCFA4C6C3759A188672EE784DE12EE81BCFCE9CBC48C7121E320D89D6BC343D5A0BC4DC642403864A14115C34973D6CA69F4CEB2625F75257BAB74723CB3B9B05A7B7FCA821E39D6935F177671F16B273BD5D99A6C72BB31F040DF4662B764F5FF05341DF3E72D35A8F26037C1D688AACBA761E9B50A7CCE93F95377F6B3BA31D54CCE4F42318E1ED3756649B77AB2F9FBD81C2AC2990346CA00C69C0A115A9A3A46CE5A3E03100BA321CA3654722B04BAFFD295836995935EA471EA2C0E04CE257ACDF16BE6047B9C38024084D6C339696D9F96640FE3AD177E68B797E66C502A5F9168493860D6C9AAF6C813977E21CB9D332D3E6D1E461A22A8321ED57AA5106FE85D79DA46878F6F68BF658DBBFF8CFAADB686F17DF942F5A4B411D780FC92762A3407F3EEBE16BB8B0632C93556846CD2A754BD9C006D39950464ABA3CDDC29F9D45D406AD660736108D0C01749F5DB083B09022ACDEDC3AFCBA9C926FA9442B4477499C0B9CECAB2B08A27383552E2952742D1720AE170938579382FD339E4CD4091EBE0E5B7584B31E58D4380F80D70F199EE751382A0F911EC275842D87F844A30A100DF66D5FF9E785C241C877F9E6C7E7A6C4BFC368C2FEABE96FB628B570C1C1F6E729955AE96690B0DA81C6438D445E29B0F8B14184EB3B5C3A3839E2ABEE0182CF5A9B4C7347C14952C9A9D973D9D1AD159E49D9EB193A36927CCABE68207F28A0F78C0B817076AA0952BF2BE57F2D62D913D75B2CF75398982B9EF4BC74D4E22AD6A8A32FA4EBE385015A18A09324B35379D7DAEC542BB5DCB1E7CAC0080A00DE4D1D8D200E726729D34363EA389ABD149415C17AC26C2D56ECCA982F578FAC9C2E6CC952F950B59CC4649FD6C4417DE6F9152E6C4C78B0B880685AB3BB83B9BFADD107501F4715EB0265A068625547D40B0C09B8AD0D69EB51C5BBF6D25D0E289151320AB4A1FC3F00802EA0D887B7E0ACDDB918FE78D98F815672B495AD9CF8B8AC71E298E64F2742AD9B17406D4BACFEC09CA3DF95CB2E16DADF791EDE16A38A189612E5C01D279EFDDA7380D1C57638FB06F8F3D00E6A365D39B9B69C448D4A5122A67DC5123647641D239DB21B6E446D52AF96CAB8124C4B990782D853D0B3DC805EC5D1B4007900E49EB2D0E10A2E983188A7BF19B0C99DCC288A93163CF5FA3B64A9B7C377213D2508E6D74574F64FF50C777FBE2338BBB2F38BF4CBC8089AE2D926217AF9E3735250D6913F37A34EB2DAD54A80276407C87C84710E0A1952FC889E6FF50723AC70E4165E048071248512A1255D555834D7A43355D2EF30DE2D799726414DCB2231D52C7A40DA99D81DA005A3014E7CE5B28395A54259E8935E6329E2DE4DBB52EE9BAB39B3839328E713E69218A5FD401F762A9236FE6F42205241BDC69E683A6897427CFE6237E13EAA6304807169D85C96BA3720A4FC7452DAA04C9C13E6DA221D5B0EE371EF13B1DDF1320E5DBD5CE3FF76E21F91121FB20F8E63399D94DA15D2BBCC6544CD1148884383D609F1AE484BC3394870002AA6AC92EE8D20D608ED4E5896AEB3028795EF2E2BCD2689C4E2F013E3992BBEC2AC936D8609EDB4288ED98DA34DC0B05AE0B60B5C19F5B8F023F934AD6FC2DB940B217437022A86754AEDD6A26D7EA43A8133A3E8A3FF56EA7F8570897AE2BC047E8043964B45165F8E6E82F3A8710147945E9A3EF0DAED0CDB15D279EF12B9F9BAF332CB480F907617ED31B353036EBE7B3EFB42F92F5F39B714278E4DAEA7C76401204304E6D45233A21D7F6CB606CECA6AE355A29DB561EBC4EF108AA029F1CB18C09A3A88FE081165FCE8C06F9CF7E7D22C3A0C46EEED41F2937AD7030976262C6F9C29FD59591DC3B787CFA5281E634035C87A7B88B8BC83C510F8F78CB91FB724251BEE38A28422B602B97C5832C2B78F6ED42B1725EE9794876FD4A935AC0F68100565F896FADD77F42252ABA83C862FBD15477029A536CFEB266A750C25FB1282CCC95FD6C5A4AA8A0D70DF83B730EFFEE8462FE9BA9690C33F1F143796097E70F28BDEDDFD4BF5BAC661319B1E654E5D5D17D578A68F28701CC50A4EC282892EB462B4E640CCD84AAE00F3FC9B0A98203B3C918E60647895F95F38919C5DC262D1CB836443096DA78E08A22DA350ACBF273EE806BD755EB9DF43EB771A6411C7D4284A3CD8E18647A2304DD8B356ACAF367925D1418CAC3FDFD45ED442B7F2A739C3B83D71A5504FE7307A37D1A88FE7CF69DF7E91F25537BA4FF89AA0295F3C47182D25AD581A889B39BBD9250D577C1A905A69D8431D11624406FC44C4011CD8C6690AAE4FF7A5AE2160CB6BBDE93C7CF0D96E0523A754806216FE43C8AFB3C838DFA975851DB350337FA7986611F003628030DF628C63DF8639E24F845174156F98B425155AA26C142BFEE5675560FEBD3519FD1680D139829394481784C435C7452E0D9AAA5BB920D83F986107868CEE2FA6BD0DDB69705D167B027BDD3C57BEC8955998AB6456BFD31B54CB548D76F9141B821F0F9156E09D128122D381A3E49A50EFD76079C119C0599B69E90141667B4B46827670253410E4C23C286D34AE7594CF3142933A4CA21B8661E1FB4DBFF18DE3771F750CF85F7275B50DD8AB6510901FF0FCCC6F26A465F4C02E899847A8B6D07880210F99CDAE037BA7F969E4A75BA945FD145763F9E3FEFAAC6A60FE6990A16EE4DF9C6B541EFB185589D5BA93FED0104A5CB8DC88618972C6137F90AF8F7999B70DF9482BD56E642835B35A8A0FAA0F9FFF1E15235AAAC3E262D4ADB8D68E37154E6155620527704866FD7B8E2D4AD99B9C8E72AB39CA71AAF68BE6BDF01D619D35747D6495A493E19270560DFA1A15AC0DD35D4F345DACF0CD82CCE1B6FD5969F957195E834C4263793AD850ED97EDAC5706236850073096BF72659E0EA637B38D412D1BD48FBA460375EFCFECE9A3335C438DEF53A9460D6B67D7C50B512026E53B9E3BF6069D622CA828CA67B89403E0B8A04B016C5FE694C9C4054DFADD69B57AEF8E8151274D74F2AF3652356DAD2FD04826757C683094B46530A5F4CD9CA7991660553E20793F480AD4361F228FC4CA04ED6C44391EE621D696B6C38EF587B3C0762C5A8A5365EF7BB03A7FC5A70FA89CD2DA491442A22E04FEDF2186246B8653CD4D10DF0CF4A00ECB9F73C5A8FDFC3AC044AC786B4B59FBA0336E226C5BA5FBD95871AE6ADC0FD1D853F42777BFA29043C8ED680D64C4BE1C6C81467D3E3849897072E99BD5FB226C8BA72526030802F620CFD6305999D59D99117CA90279BC39B97A1AAA5206BB82EA39148C5C7F60E20EB6516604224A71E579E5F848751FE2E85FD51B9D5F499D3705320917D7DCEB2A1C82C9395523AAF807363E7FB65E34C5FD3550336D5718A0E3C5C5D52AB3A282081FC5DC30CBFCF1EED0D0397EE4AB4938B3A7E4D5DD088E88CED03A73BCDBE9D75E7102AD4E18EB565290E35358798DB9A1D1A019C2155FEF3D02AE6D7B23041CFFFB97F9C98E62003564ECED8807E521F317600FEC9FDAA88B59B9B7BC74DDAC0168EA90F868FFDC00D657BD4EF4BB415A90E6560762854B67A0577E11AA6B8F66D5B44845BC108447E54CF695A088E53D5AF8AA53B797013267A02F3F31691F7497C31E1FEBD573A25F20CEED1789D84084110B65AAF7F709D6B5D95B519737E213DC5FF810C4BD968412C3928A1388D473587E0686C0F5B795C3B7BBFF01566E80838D3DF2FEFA384628242A16B73ED558A6FF3D050809979EFE361C0690A101E40086228BE2301867CFB425E1A1011FFCCD4041AC2CF57254028A3EBFDBBE5E52BA19394895B89A6F7C24D14580D8A883E6A95D7BC957FB860B2CE34FA1D011BE071B6DD0B6428D74D90235899AFC827823691305F54023FB37F49CBA642600E014C751C39B46A82B3FD106AB6AD55C166309D7FE259419E942823027A5F635322D46324F1FED840FF20D8024A82231683CCB83DB10AE9D805944D95BFEF8920478891FCC66E82B4DCAD933622A0CF1984C891CE2F37CAE4C485F261489DF023F768242C12482CAB4A3B92F233372C1D41C3E142456D0E85DE560D08B0B6EB74BE5014B944FF199B05BEFC74AE150457E41E01B50DFEF2C7861D401F77EDF17E7CEE6FAAC0E55586B67260A8CBBA3CEFE1425639336CACEFCA60305E77D00F2805F71FE72568288426F02DB6A162A26C6AE90927970DE83F1F570EE758161FC5688F48CE72F84AA71CEDCA1CBBFCA02A1B1396925ADDCF81E76C2CC7EBA82C8A5B013B8324CE08989C85555E378DBB27E4FEA5BC56801282B493D09895E588FBC65C101FA4736D96FE6496001684E59D28BE1C4DA0A566FFDED0A22DFA4738C3B47F1F45B92BEC7E80F7BDCE914DBB2F3D806BE027F9396F3DE4DA2D965D388A5E47E01E8D597D58E8C0EADB05A0F5440E77C76F83A035142ED6F57343EED40C16A9F3FA48996B9872B8240BEED8FFFB8B2B751C6FB27505F0F30223CD6BFC04F4BA5F259940C48A1224AE4D57DF802ADB2FDB8C196459601A56F71A61D79637C920A9F4E1740234ED60693AC8CC75B1FD5ECD164173204B75CAD248125DB9CE3384D1EFF2DF913682F957AF7D6B8C970669BB469F9FBF679123A577B2A41566F017CC9D49BF9C00E92FCCF10B0C3C195E00146A13BFE058DE39D855658C6666383F74673350C93DA68B350F5B6EC9423D22798BC7C7F48E2B71EC333517DD2C708789F4755F68986358051B76939ABBDB534C7DB0ABD5F017B4A9307A46D82B6CACC285464D38EE77808BDD83684F85006E05C779930D3FCF08095C9339F98C4E674444C9EA2C8E6E2C863DF6F42E7E7D6730FC8D9B7767CA2C40E9323F5FFA479C126DDCB8541C750F2F49EAEAB0139B7F8A9A1754DE41247EB2488C2638020BDF727B040CEF86EADE4BBB721C26383185CE0C9A14F50D1E293D8B5EC03E81250D926CCCBD5BC53195A7D20994EA952A0C4617D065A8E64D8F15C187E37DB8D858FF68FAA8B04FFA0CC8354F8ED867B23DA10FA39D0324B6BF131E5713B96834D5A7FBEA02E53FBBC26E334B1C5FEDC7B385319A6F91737273143B00C786DC8C27474A4C64B00A512C1EF5DECF4DDF16F0147CB60F7AE07E68E24B589FB573070EB149858ADD70D9CE6B054B9B3E027291B1C538C67ED3DEC48A1A7DE4CEE827DDB3A913A005A9EFD08B4758DBB99B4FCD248883C8D0E2A03263B751A86B41A86214D79652D013EF903047BC08606013111244D6D03ADEFC5B8AB5E84EC348D59D353FC3EFE28749F8D5BEB99B281A1756EF5C6A40CCD04416AAE316A1205A0062A864FAD195382E80DC617D65125129F928DDABD45FFE31709930C01AC3FC6471F999DDB08F4F40D2176EAB177FD10A3E2133E2FA584C69DA125F420047955D2A1BEEEE39BBEEF8CD7BE057BE22D5B4979A8E065E3A7540384E1163AD20E18EFA547D26E44145A8792E3CCC0B6B042A9AD73B39C8EAF66E6CC1D77802FA8AAECACD1EB3B6B6D7254A54D8D85F12CBC8047266C5CD61C95BD3BBA344A37F482E470081727FE5D65321A6B1148DB77DE34121877F79C94F7331E1EB7FDD536177BAFA818AD9844A12F793A4402A8402F3D4908F96360A82EC8430DDAFE325EEBCD40B47EBE33666B34707C5B90AF1059B0565B6C9F91318F28535D837E29E088E53C39038BCEAC69BBB5214DDA50E593E6048E8697F4A1E5461CA31BAB28C949DE4895499B135BCF57150278B084C6DEDADF9F6E9706E5F89A65791FCB897601985968D0BF4DFA454F9BC9C5AD8755026A80FEA0DA6D82BA3BD72AF0C12C6EE1C08278661C8EC886CFC6B2B5CE683C36B5DC71117CA533920E691718AB5015E7BE083BABBF3F21E510D681096B136BFA3EF9D9D87A0AC6C0A21F6423E2DE0600F000976B31AB1C87D62C99EA920CF80B0DF7EE40421B7DD1AA10385654A04B5C9D8E45A2396421A91554FEBEDBDAD8DE9623BF7553B06CFB764F551838563935AC5F7556992768C2AD57BEC47D1857B0E8750F5DCE9BF2825E199256C161C70CE8F65FA604B4AE8F797BFC7B9C1DA00802CC6904A3C7A0B630733DCE8CC1669827F07C3707E79BA059CCD3A8681B3E1ED44218D1B0557722CBE0219EFDD29287CCDCBF62CE7FE233A882E76D2B047D5975E0032B790CA01C55CD6EA175343A3B969E5073863B22BE6BDA32AA54F8019B89D9FDA2D4C97995A327CD3836B03A1C3CFF3C59229385AB7E26C47146DDEF87F3737B0845F7A610724631AA3D53D833084BEFF5B76A3F3E4445569D98E5F9863372F7867BA0137EF59B6EB87D4B0F1736889B3F253BDEA23D7E713855FBD2F4B69C90C4EAB271F68860025335CADFA1D66B1B15DF08FDDBFD6980545D675BF6E205AB298E829FC75DC701DBA0707EE502A240E208DC22CF38FC76A0D625AA3DCCEDD55DD6C28F83CF2FFF02CF8414BC153835DA9ADCEFC77BBE87DD8C3E48747ABCBD2DD1F0BEF11A73CC5C21B054DE3F68B070AB634CAD123E1D59082B66C67D69ABB3BA89CFB5DD14597A6612F18FB372535EE384F28DF5EEFE73A7560D7419DA48F176F67529220E5C0851E5A525B219B05AD08D25F0D880D193A49081440F189D16B57CAF8668BC7B74DA4EC6C9DEDBA1CAB708492C295B481C13428914ED246B3E670259E3FFBB446A6488CA3B8ADF32118D14BA578215E25158A00014D9CA3D6551D43C3ED9565005DB17F16F8CAF4A45CB48B9E615C8A247D41A77B354F54A9F206EB475ECB7C69905B11E17555FF9148FDB72E7B21F65BA7BAE296FD518628390CDD1C02EAD988E24AF18093F905BBC2C25BE559D5606488E6DE8F59C72E98CE38139F33732F9C95B827FB0E98B0C91D6424CFE11113F69F44D0A79821E15FE2DA83F8557BBD454A95DE9C689AE47CEFE1E85DF3478B713CDAA5CB6457079493E240D85A40BA7450A7459DD2D0E713F6061968D184561A4CF121C19DF0307AB0F26A65A4E09F2D46A9A824F085F02519F668FB334501BFBE77FEB4D3B482879AF768666C5259DA3510D06EE0649C6C1F1F3ECC7662A42681001FCE54C42676B3E8222FF698BC8B54F1A886E4EB6C4A1B57038BCECAE40E68F5CB9C81B5C2F2CFD8A829DABCADDD4C06FD3FE38F5482EB82FD870A1674D6921BAEF153FD63403510C00B94F0A214AEDE5D68FA4957171E6CF5658FD0AD5A4C74594364015EAC56DF6307D936A02CCFFFD2F3CD5E082EC266A8BFFB6C281F2391164263A6E1B4A083F189FB19E5A8C2C6B6B8BB02B50D336EBAF3AC726995F118A4889201552A83CD42D8F682733C8633D37A3591675BC138EDA88BE56B0DC1A5355A594EB6D63309F09FA4BB8DF28C2C9F7BF8FD4C2F3DF98086E840B376AAE9B47572CD1E281FFF714B722D68F7E7C465E217213745CFF5217769EB43D0784172ABD19B9CAB096F8A88C0316CECA80C13141FB7EE47A31795C6AF41132694AA9268015E639B30D19F0B7AE402C8D66C404B4C0FC8F48EC59503C17FFDDB5AB3C2904CA8C7F904E07F1A31042E379E0F97A728BABB1F231558CE34A0B68767A2A488359D098BAEDCD67D0735B1C01725EAF866A24DFB9DC68101DFCF55BDAE5B721CC0D4B63478B462EAA6A169621BF5997F30FEB86733405BD688195E3224F784866729D45E5D7560EB889A9422E758BD410E7F232812F01AD0901A700DDB38E4B87CA02895B3CD2DF1E12D78955EA3F31B985920D4B19389B8A83D3D5228A447477A99636EB2534937C2B3D49A22008A1A0013A29D39F8839CE5BC47D970D57B5923B5003DFF11296C438B87402E93F410387F55449653D3E437F5771D2F41808E74A39F92FCB4C5F1AF80EDE76908F9B20CEB33C422AA3520A7F3486747C10233B3724E1978086752FD78C3E0BC6457E311FAFFFC074EA5BDB7B5D73A3E1DB881E7486B8803DF0D30ABFF855BE06D77822784692182B69560B8CA5EB73E0559DF8D4F58FA697533F1A7581D07D6A43A4FD4A3062FD38EB7070BFEDA3AC23B570A0A2228CC7F21BD9B17EC2BCE6B17836B8ED8DB599D89BB6F587DEBBBB42E224EA8AFA74DECFB309395A65E1CAB0D07E6E6BA331B1A639A29C5BB92B61294DAA7F030C51398BA4927C1FBA94009735BBADAFECD71B31FDB511BF41F1DA43182FF7359DBFD6B374148D97A04131C240ECDEB4649658347348142DD584F1E3CC10C1764BBB3BB86E6BE00F04D614246A90A1AD466FA9D4E7A45B375829874A9EAE8CFAF797AA3F74070C3356A9CC904726E0CE67EFABDDF48AD54C6C6AB8D7F9881B5D1744AAE1E00DA9AC0ED939438CFB0D61CAF0DBA07386F6B92DFBECA264716701741076A56F9677819553F011DAD0C517D59E573A8AC956D1DEC2953A54E0166BD3402CB17C46489074780EC923DAA3F36C99C38AD893B84ECBADA910823E045B4D3303F46DCE53D34CD3C85889FCDA5F3ECAB6182CEC5B45B00C62F8CB034B507BC1013B6511E1221B909DE20493EAAB148176C4A131EBF209F33EC88AE0DC7C0FD2F740E565FB9969780AAA15DCCEF13C522C82B4BBB7F30CDBCA19CDC39E98B48603D52DFCAC7EAEA7ACBCB5031666259B03FE98712E6CF03A55ABA84ADB668541849B5F7EC6A94483D3A8C377A5F49169408327BD8E6529501388078582038FAC6E72986FF98AE88E1EEE0292CF253C134087823FC9459F53B502490E086E23550124CBAA46E6396209E43E0402557CF30491A0C7AC48B9D132DF743FEC2904A507886B20CDB93453621A99AC215BCD7748E1C9B13E411569242413072B41820DD089A4CF10C7B1682A77E176EC3C2E6604FE8D44B80ABCEC857B2AAD8231C14EB13F2A5448E916A9F435763894E1931C95F98CE33C166AB993A664115509A5E5717A1429D0EBFD52F8B36DA3AE33AE38BA962338C430B909247332EED2B299982CC376D9333F15016E66E36C118251B34299E3A650B74D3A3248109D7B84B82D6BF79FBF6322368AB39B816088110691309B554B770757F32EAA60FB4596710BE3F9B966A2F398C05D6BDB55BAA26D9AEFBA9352436F59BB5DDF284A0CF8364882B2B099D7CA2C42A98173672C9EFE25A84C5B284F8B8EE23200DCB260C38D3B586C8BBBB5C21F8EF91040DF280B042E6899027F3418A9BD04B2238BDD93AB8DE02335FCD9F531C48BE13188A9A0AE4B0C2850D222568CF066718FB89E9EC48ACFF73A1E2B39A6D1357D824929BD156480A0487856FF5BD6E842A576430B2EA903EEF20A7E63DB04DA5C33FAAF9A1094E5FF131FCA54394F626059419AAAA225D0AD613C98A0A694302BC73A18EDFFCB77E1043FEAA67F7DD3D19C108B99BB00FF1E88508BC2BDD4E7296073C10DF2BDF16A270E363943CFB98A9F6DC06A31BC3BC1C815B2CBD4AA3F6912CB37E8DFE8EAC4425DBCC840A8E9A8E15C34CD17FB38A1B7F527C85A69F9014947C91E17951BED8DFD675CD871E46D0737AC69F90E64F288C9C473D92703CEB1174DF817879C7D54C4DF99C7D1B281197946625341A6689D876B7ACE62546FB473722F3E93B9D9B10549C65A7C6368DECAA18C3595223AA65C547BB26D47173C958565B267FA2F73A3E743786A5FC35C7651E460B48918C1AF818D624670E6A7B9279979EA65C94108B17704C0865CF2D47FC9C8DA72A797DB97625A7285C4A2227E20FDC7E36028B3A25D5B23D391B6EECDF0E126E21965CD24E255470121969E9424A3E341737ABA623BDB480F68B61E153176608FE320A711324339121B2B4C8461FB4FFE3D6F77E93803EBAE38B752F12EFB1C9289142D5F713F0731E731404ED1775FFA435AE672CCA0339D4ED2365B03F96E49EE8AAA32E417CA49B05C3862077CA3E06E585B0CEC92AA555EDA01E5F53F9458236557EFB8408F989F418C236C576E12A1843D31FBE4E68FE4C57FCFD81707C9F86C8088AF28A43FB27FE7FF42F4582A608B4D27E4D04BE7939ABE53772EFA47C88BFA8792C5AE178CB21FAB664087B5B7786022498FFF402E3E1DB5A61AB1BB14E10A6226CC3264BA58C67AEE884939A6263981F31B870E92C32DB709BFC90667DA06F6AA522F0628D9E91D3BF4CFDAC3ED78ADDF63277A4073C69B4E2A01005C54649DD69F399A3A2971C47120E41C0816AB42B16F18EEDD892C235017DDD490BADE664A46B96F87E391E5321EC885AE82215A273A8864A3EAC35962A7E7DBA2A2BCE1BD20D9E5D7BD32D4A3CB94BE6C6975D5C68597026996B7EC5F1BD998348A5F06A3BE5B5FF3FF5C9C02D032F080BD422C7C328EC5AE4518A8A58A9916D419EC959A7323B1A04E093D991031F33F9287AA8A0F7FB720703CC1CC4D3C751C07EB65B2B744431C01FDD1F0D3127405EC64C81C8F6E6A8D1874CC83798622CD759D2BFB509134C7017EBCA7AD92BB9563049B147374D90CCDD6D1D4F6ED482058FBADD4B395642B0C5526BD837B4D10E776F1B4A0C0F595187B7FA51ACA303AC7165956036711969FED6F53E6DCAE39188B8FD7D55FE69F7D20FB1BE970E7F502B1E14E9125C2EEC63F6CE140CD0913F79AC9702EBB30117CD55609F32E7BABF4A6600568AF47D113CB1FE28AE03B2829486A1420E67F92494B896AC29C040A9BF139CB3AE003D625359E552F9710412D80BCB7C1C2811A8BD964150A806A22B6E59C99CEF82011EDE90E2FBEAAB9B98DBDD8487160202D9697E31FBDA589488E31444B251DBA9338FB90A91161CD55688B971E71BF00364F7FC566B7ECBA442B4F8A5E6003BF56480E3D386E96B9E928B5E5BF25960CE55652D109952245FE05CE83F54C311D3E269E3A53BBF3C1DF86D266898BDC8DDBC2D86EF7A9BD81F2FA8AB51BAEC8F779094B814903F818FB3F03E39A6E4C9AFEB86B56A6727D07F8193547FBEDF34A77E1B272FD29C63359F8B27B22840B6023649A65CE51CA2374CF20D11274166E4202C3D0D889DCE5C3E46E12205025B42608F10EEF5A4A8F1F2B2A21954C0AEDA542A4FD44DAB0E4AD69BD253345828CC1B81EC745D6156C035A08BD5428296C4CA628526685CA147707E069329CB278419398BA168D0209F6674AE9F747ACDE498E7094DA29EBB4CBEE613D8398ABD1C262CBA4088872CC1A04645F6C6B26838695DD8389876D044792099E483B741572C8EFCD118FEB27B3F9CD88E9A3FA0296797B18E17C62049A8A027E2E2E1930D486BCB7979AE8DD7580FAB1C94828ADF3EAD36D2A02EBC1D80C6346B87733E30CA944F6A11FC95361B7A4B63A5B5B3DA88741E97718E08B260C409078E8388FF57B7DCE79C68788B8A7FDB0A8DCA8119548B1B0FA2B6DEFBEAEB43866802DD2B8068EFBD00040E099613474F4CA7288055614BCCC4611A61BBC049A5CF476DFA53592984916AC71F946599896D613468E889B8BC65B3752F05F0F96351ADB20060225CCA3CF061197278BA8D2EF427D6CDF0EB0C1E6564522BF9B2ED12120EF55825F5518E37E4758C2911C48DD6F3664A63728DD2F3A13117EAD500B469FD9A522328D196FC221228308246CF83EB7E094A688A626C1E26B4AF3C47CE9D8DE2AC380E68F723B193230D0EA5CED81B54C26E7D774CF8E54A610D48DBDDB43584571B49C315300DBEEA8B26EF96AF11CEE0E6F2AD2D9A72469CB6F31633E767222E1FD9171B2671900A000BA1355AAED1BFEFDDC84C84A5FBBE20631EB9E5AAF2AE64506A8A3E31C80DAC27D9B756B144420D5576219BFC3431DA6CF1469BB0E49FA301486F03B28A86F7704C8D05303BD0CC6E33BBD122BF70C3E51F7E7B5BF1A0055D2BA6F33D75637AF70EC4FF1C825149E72F88D15800A5BCD6A0FC8A398D57B3E47594624684BD17361FF7595B606147E5357730645C2574A890047F762A0DED98279706D7516A20E59AC41F21CDD25963A6BC7445228348F473A81C5CE53A82DB0CBD842A25046D58982090B5527F84DD19F476EFD98658728A223CDEC2F73AEDFD4B9032F888A9F6722E0ADD748987AC762D28EBBACE5762B3AF1F30E8B8AA200FB7399EA7CB97470C8F3029F21AD44D5247E9DCBF01E2C0A3BFB30CE0CBD72CEBC4A59CD00152E734AE0A4CCC1435FB469B98AD3556BB3EBFAEB83F70AAD5BD7757A561CF11411BA35D6DB1F4FF6887591E4036F8A65C33F3E29927E91A6C3B37E61A1D8C1AB72F93B9A6CCE40D2849EFA553EBD8DCE610D101B1FA66C0E58D16FD192795072B68D513EDB4158F2628C1F8DD6F27B718FD4D9D853B5CBBAC931755BA5B44BC6898A27922DF2D21B3F12DCC68149D8613CF6BC0F2C7A86FB386DB127ACCF912DE879B99062A4C5A40C9CBBBBB0780C920217EEF619C0B3B4A0568F10ECBE8135AB42DBE77643BB5896F9A6503D34FDBBB7094DD1EEDE79ADB450B4B9CF23149918986E7F581AB799DA2AFF24668E966515F12EE3D048B1CBACE339188C1E927EABE5CCEF78948E389B98043774DA5122336403754710B'
		},
		SiggenCaseItem{
			tcid:      6
			deferred:  false
			sk:        'A37C1089E319A6AA532A1804941E6BDD41A2D7689B0BCE347B90DAB5EDC2519FB44879BCD2057FB09DA59022D12DA09B9A86442911A224C58C4CC574D089A2C3'
			pk:        'B44879BCD2057FB09DA59022D12DA09B9A86442911A224C58C4CC574D089A2C3'
			message:   '1DAD1F2BD3EA2108A1B6D7ADF82E58ADF660695E15E33F17F2AA42352005875607CCA09CAD1CA75F00A210A84106BF996498376A0B94C3BE49CC477A4922AAB25E19B3B8C8BC452ECB75F3D9A189E33A248B58CBB7E670BB846858F24A72D5F47BB2312540E425BC64EF517C504826A2BF92ED1E162664903FF49CED78A91D1DF24321C82BA2CC12AA6EF21C77AFB02156D09C678FC7379D7A5DC80DF6D02B560BC92B00697D725BFA7DE54EC3DEEE070193BDA30028E61E438B459EFEC78F90BCB6FB66B7B1B514739D9076E57B28BFFCC7D48660E70C062FE3B11E91E6F98BF3CBC9EC9EEACFD51A1E8B0D2F1501F5AAD684F752835B86A29A518686CF32FEAABF8BE670D29681BF260ABB6DAFA0806938EEC3E5A34B7FB139BE356C8EFB25D9F9BCCF956B2E989A6A9B9D030DBF60CFBD1582F40BF7668F21529E6B31EB5BC30DC82D0F703D7FBBE3CFDD0ADAA103D8296657E9BF33A127CC40D3EAE97C6A47A678A410988A3615FF4228AD1E33D0F53C88E79B32013BB2D9C69AA6527EFE0B7DFC3DAB97406111028AEBFBE67BED66E72668E888E743E4233B51F99C389FEA3E0E280C99B71CA571708276E65FEE2AC036DFF2683C1AA608D762B3E6D2818401D15AD4A5AD9CC619D125A28D4CBB85EF37CC1EBDA0BC99E3CEBA367E357796130FC2A2E4DD618D549D9325D6FD74C30EE0E85D699594C3733FB2073AF164ACF7FB9F010FCA66D79435B3526430D995D5F528E2E16E92B211D26C4BB4F6C207EFF855AF924AB836C2C9CCFB47A696DF8B67FDFDF954A44CAB324CC70029A06130FBF8FA0F64FDD3F3213685BB3DE55D996C745557F302E8F36514901EAB57F94F87382D032F4CFFBD55F1FB3C97B1BFC26A725722F0E86928FC2A5C63BA29E41D731D6CFCA8C80CC49645405D2BE41DC1774A4790746C6CF434D5CC3C109602954E2720B572370DB203CC8F5CDD9EFEC8676CF9BDBE334493D2DF33B57A0F9026A21DFB29AC842D710706C3B9003FD4688B474CA1BCA5B34A50CD3AA0A814B8C6858F9CB106890FB30DB562727D95610C80DCCA33D616B53ECF02B2BC383B276A78414E614C5444557A22B771E4824C038A72DBCF7F3107D4F1E8064BDE8AD5C52747F5CA99EB7E5CAC4964DDEBA627D64D91470E004FB16D0BE74DCBB1F09FDF00A3180B599995D180DC1F319E12BC3EB3B73C7E69D66840534E632EBDFF39CB7A03F0A7E5DA8E8910B1E4698F04BB6F160ACAEABB1AE2F04AFEE6E723A5826446AE355A81D2487DA2F8984CC6B33E393587D43F647F79B05E72792E583081A8FDAA1CCD3EF1F6EA492E6935CB4062C42C3F18A54E7F0F627C744C78BD92AC0B2D638D29776A784D2C23BF73E2F625AAEA37C0053CAF0C8AD39338B63F230D09A24B2BF0EB4CFBEC4454545B0AE3F6B52B8C9BCB9B4F57595478757357BDA2817EC956D8AB503686025C549408600249078F73E2A48CD2F924D74022D3FE4898E85DBC0C2CFD449F6E40576E487B30959A49719F558BDE3AD683D6F0EFA5C75ACA9C0F39F69D92782FC96D83C6A97CFAC730C79A581335F897B2A9BF767469DCC41E18C576F8C562E3C9B38B8376EC80434C6458818B78E3618632BCFF7541E255F1FAB32ABF472C894925D0F6977FC96EA935B757BECDBED14285BD244FAB099AA923023F5B297804BC174F4A4A25E744560BAA7FDC8C78F4390E54384BE8A098701B1C7EC31F7953B494E337C1F8DF96BD090DF04479B5C5A2C65FD47D2C989F4E10432ABCA44D63FBEEF892511ABA98E3D165E487EFA9B345D82310837542AD2634527B91C36822ED94E0ED2DFB9EC5D6E24ABFD9BFD4A18CD4ED24C73BF8DBDC268DEFE0907B2D913FA45B91358832FDEA4B7C511ED3B424320C0DF0F96192F07123B62D9BAF225F9BDEAD74F8D399E2DD1E28CDE94CFFDCBA8B90B3DAC86FEC185465CE6A0F1B1319659D1DB06FAFC2BFE8B9684EAA44D6F2203DB7C33BC439FB5EE3A89659CA978677772E23F1FDF84253EF9F026A4BFBFCFB2734A7A28A9193C10FAE67F216AF87BBD39AA641D21A55E4594DCC57FA0B0D4A9AAD08525259111E6FF50B53DC9CA1BBF7FC76584696A93086F9FB9BAF02B61B02438EB76B7EB849F3EDD87B4ADCDE55E97C5AB1270F8E286573D00BA3040B47715630BAF18B3851AD9D68D4BF0EA357059FA0BB4A277132FE8043A3D066E75BC2978AED34E3F48A37A4D898428DA8A816A0728A60CDDFFB44649EE61570F58636AB6268B7BAF8772A00892922B5979D665814C5EC1D06240041A82C5B1E8AC1CDFB4ED92A0F012B665FA866F1DF3CEC91FA059F31C38185848C78B8E55ED6D2677B085EA228976BF845886EA28BB078F98D8B32F1F13CD55AF102C27AFA70EFCD4BF2A257357A1D2CF6916E98DB76874FF3B2564DA41D591D60941C46C4628AB4214A1812006BACE4D9D60E4A5A36EE0D4887DD842510176405A2C3E25EF60305DCC8CFCA83D0D6D0377B5EBB815EC023777B3CC767667CF0149CE2D63BE45F389290A81B596688854E44EAA1012C00E779FEC6BE2E959684E328300C552514221D60E882463A213E396B5CFDEB601945A838FB50067D987A13EF557BA4C1F0AB42D6021A72A920754ECD3BC710A97339A3D5CE46D057F81F7A5A2B66AF700B74326DA75F99BC1B767ECCA8FF9C13D53F5505ECAF362318EA359CD78D209E41F7CCD7DAE5E8C93E8F84046AE9412EBB52E84C05F067D74C0D538F28D84CA07BE8B5E92D5765BD8B5AF6538783316C795E74242D9C87F7E0F92F40A3732335E30C889B55BB8C307715E88CE748D17C4DF6034C0D30AC04840BA5BA87DDD274E6DE9C58FF7F627DAA8255D9A00B0286B4B71D76E80A138064881AB83937B3CCEE8998EACE85336B6DEB5721B1118C9EC3DEF13AA9C1FD7FC86BDE32EAD06901A406EA2DAAC564A5F1C638E689DBEB43BB0588A23857D2D9B742AF322A2532A5D2E1FC9C5447A34B8029917C9BB5C2779E09581C753BE2A0A33E754E11E4CE8342D49B4B53894C1321FEDD1BF776182C91C117F9A975796D2C5026A05AC5495E4589F2B4E15339B6020191EFA80FF0CADFCF145B43140D35887C9F8C404F14B3ED862AE840F8FCA51C5B0DB6AA02E9CCDC67EF6E7937E5707232ACDDF8551110B73CF192DBCD31CF3E8D9228848067345A98E15160CCEFDF1906B671C73A33AE84923611364364BEB84F3B6916FE7628A374182C0496A2EE4D28D6408BEA1F79F6A827FBA80BA872C4E5E802BA3D07EF46415BE7B42A57AB8DDF1DDFB628A4A152F5A61DEDBD6AFF5BCD565B4230CE6B078C682F8B726F9DC614B8130A033F1A412A3389A80F7BAF71E65924C71EC046F227E3F643E5CB867F4F2D696DDCE6B4F11D7A0276C093EB82AC1556F8EEEDF47D26EFF0B83138BB2DA94A3CFAFE5C873D5213B4123E6CE2189C287BA1F82FC98B2767C963230605D28D41E2A3AB87AA28B74F27B7791BE5EF5314BF360A486E8BEDE781A9843E8C79CB2D2E245C352D5B5E86EA67BBB673A9114DA2B080D000BB653ED8D9E209AEA1B6E36EECC4F63DF6C440060B04D4CAC6C164B333E0435D391AF31B992BF29C6591EE3B857C340DC48083F3DD091BAF81D804CB7E6F4090F168EA21D2BBBE79B81E1026B355A2CA8CE322737034C5243CC6D658A4AABA76B8A2912847C1F1E7F4F328A32E57755730A97539E5F833829031E3C3A2B36DE0C23E7D28ADD274021C086CA3B756561F89790B128B7CB536CB3EFABBC40EF06197E0FA8477FED13BBB01B69B2FFEC18BEDA7D1921504C1BDC3F5277E0E2F03D3A39BA279E243C75B0B20164C39782BF2BD08EAC8E193FD3959DDC73F5ADD5BD24DEF135AF17E94D76FB226123E1A9A8A34815B690251C3B6F693F8761B370E32335567D3025F741872EC19A44AF4CD5153E376680F8E27B5C315BA659706C4895771060B6CED6DAAEA6BF8290686CCB0F98F7DE0C065A33961D3C1700A5E846B16202B17A5C6E1D0C337CDB3C889898586C5C41B72DBAA8288ABD24DBE31E1B71EC1B38F0C5376BEABEFBB6BE72CE5332180A1EC16A22DC9B0376B1B848CC07FA2B4E0AEBDAA0528B2DBBE9FA55BB9F4C757DA7FB0836CFE70703A127C2899698F61C6A121AC8BFBFF527083A19D39EB49E7431EF550E06856015B48A6057A225E603DDF4603DB0A75CFCF90ECC200CBB8E117F74BF8C9CD400CA4FCB700CBCFE25C45A169F1CC61DE8E16BF1D2074FAFE124872D45D7FA402A7D11364BA998C8EEDB160BDFEDE0053EB54CA9DCB74112009B7508C5ABC93BD03A048F2204C3359B38A92329404B563D5CC90F13DA8A2EFC334B1EEF340197FE3F5C2B442D6207C4508456D64D554BBA643CD743C76B3C5548AC841C87961F9F8F707E9BF5CA7A241CC68F06DF67A8C757A6854391177EADE8110E9786248ADF8B264DE61CA350E980686B3619247647441A311275AAC5CD669B3F56A40A9C780C982B55BEECD198C8FAFE56E4D5492777B292129C8777B68BFCD2FE3C29D47ECF400B524BFDF9E63CDDA9FD5141BA39897B7088795BB807FA7743B8C30E6662E84F98AF0EC292F83B1B7E549F722DCFA5960CA28CCCCE67EF1A24EEE634F1AB22496F8F016FDF861E0D5547B3A7221F5629FDC4B998AC57DEAA1EDE58B0F59063220BB19183F9935AB63B3914AD020DF88DAFEBC554DD2DFAF1130B032A4C593669E4C5B51A9D0605B31986B6A748E1A51208A51A3BFA47E7B0CC3E8A0F56744CF1D06D8EB72FF122BA17CFACB4EEC72F9D0A69AE894B16C7737CD50BCFC02D82C64B956E688EBF8BA73E6542C1CB6485D7FE4A2CE93A88974EC61D66ABA8512F6A91681964AF1DE73742D911E2559D80E370A420EF98242E650A1D8665E6DE804047A86F4C48068C1F39C50D68ED915C5C835D7A28A1671300A4616B2B3D10FC5041FF73B1FA0430FADCC246AB24D2C67538B386D33EC23FCB6A694088F168D17060324BB40695100A30A8FAE1227D79F4FA6C941E915C928DA38A471A1E71A3C7A379289ED7C0D1CCD2283FC15FE355B1736F0AA53084F988D11374E861E232707A4AC4782EED63F501C4939AE563912872B90C40E21E1277F1578C3BC5E39165B32524E10BC86A7FAFECB342FCFAD05D5F4ACBF357F5959F3BD040996D03E1C5079085C5B0F0633EAC543687BD4E4841E0F94FB7A8990648EAE5E17F0706D3E6646091453CC1469EF2648C5E4E80751D4F479040FA562598E5C287079F55A338B28508226B9799713A3A0DDE31EC1B71FD70C4BA3F966B7C92FCECC64270D8F032CE4A5A02629E13F1DFD765D2C895C298C9887855E5F6FCEF1A94F9AB9B5101AFE096C7AEB44B75E92A9036934A8737E69851938278E0D985E91E4DE8773E92066AA069F08C5AFA6D1AE136BF8CE5FD588D70EA2D676C404A974409AEA880DA515FB38937EFC567728EFAFEC92B70D9E2BCE679519FE1C9E3E849B5E3DD795809BA622056D8AA3F06D28A1F215038945D37D728009A94C3801A51E21ECC39FC9E2C4F01CFCE01C9D4E713E66371D445DA68822DDA178448BC21FE68928F261AC8ED81059612FCDF55A13F84E350F57E72F47144D6F2EA2F31E514CCAD676B147BF73758F0574A5BBD6920B436B62DD0FE9BC00DA39201F046816CD06EAA488655764B1121E41A430214E6E8F320A09EB57376E5EDC08AB708694D1A9A4C70945223E4E754E3446581ADCE2E591A59839C071CDF4E9AAA4A5D9FF46649ABF0C04330035CB43C95D252B570880AE8570CCF96B69B0CB3C455809923EAB5971B0235D906A017291A4292299302F02AD3718ABA0D64AE269959E02A85CE8F27FBE5B860A2EE59E1B6DCFB54B1A61DA4800667A312B17CD372E8B76091DE0615A753DFA0B770213B14AD6B8A38110F40BA71F88BE4267BCB867FE0D4297E8F22573375C0F6C82678924BD99E7D034353BCD0DF10F06D492D14C678DDF8C386FE3BE88D8B74CC219982F8F92D439091FF5DD9A7A06CCB0AE4BEEA9D1861B9718B692D3F1EF2A12D64714BDC0B520807B1EEDA976A5EF01B6AF7802C923092D56EF44B355B5270C9E533F69078260274EB8CCDBB371865D6AE78818FCC86616B11C4020DD6F3948F9A01AFD0359E83FC875CB2F39BB49961021228FFD21ADB85042C3F0C2299D1AE80696FD07977F8C76863AAA81B659740C024A7A89224E909E229482E65FC5031F4DE6922F56985A9CACB14CB14CDBE5C5A950872CBC67CF98C654A0F21B3928D2ECF65C9C1E1E5D897737F1F1E756F3C2879D1F8897EF16AA83B04DB422D1D39DA233083F9E6D62C8D81F1CD31152481309C3C4EED6CB05F535FB0980E636A9930A02442F6AFC864C8CF5539DE44BA58D3134EBCB65DDA0E763733B24B9EEBE2CBC011FB7DF7948F48F2ACC76B26868711FC36FA563659429BA24A9B3F01576586C06064DBDC550A0DA4E31FA075A0B0C262C3A2F462B32C24EDC7C2F1A2242C024D3D1BE758E9D5AF2B6D19628E3053654C4D533D69A2C3EC47BDC5B1F4256ABE459DD0D905FD1FC5F10C97269F73E2A379C7271CE271A02E0621E468AFD6BBC293B8D670E3DD2C635A45BF19C0CA0E2C267598BFE7FE772C1EC4A632606A1BB02667F0ADA0191902771F1B699DBEE2BC5444D2CB86D22A9456768A0CEF938265BF4CC8B386627109311F821292DD9298C195D5E2CFCAFCFF1B870011125A21F921AE373057B4523A37A28683C1461B6687AC57119CB403F67D2067E89CA8ABB7A35368AE342A4528B77296D3B17A1F836F9CB9CE01D54C9A4C7B5AACDD09ACCE76380DE0D98B03417A68E6E94E5061D7CD44E2397721FFA1343239377BBF81AE5BD5241341ECC851D620E0018680CC85B2C66C5EA808A3AA5B4FCD91DCD9726A6A7D6A1AD6149E29939A321ACC5AF0F1D41600EE29EC1BC5E00A37E0066BFC084BBC5C8772A09BC3B4864AC3CE93A4933FC40DD8D1CE16C6F4ECBB61D842AFEE5E00AE70EE30B5E1EEE2AC30A300A2AB6C0032B65A5A08FA3D4AB838827AA650B6FDD4713F1093628A5822EAB85401AD153DEC8EA366DC2271ED9181A3303A01DD6494B4BDC7D9589EE61D268C8AE7DECC5B78CC8C83C55BA2824918793258978EAF759022CE088DFA690278C28EB4BAF60AB3FBD7C8B14304C782B655D3B1915EEFB53145DDE9805750853DD6CA1325489EEC2AD3A78733E0BB7E1C5E5FEE8FA6E942E5B3FD59E23587A36F0C920E72D3D1163463588A91C5693E9FC01F07FABF81DFE54CF7065EC35F835E494C9D1F5B4E2B565A9E1176CE8FDCBA4C1D31B8D5ECAB99A159C10F3760C274DF492192137ABD01D7EDE75B2B813F0DF63DBF95C462976ADEB08A0840034431E93CF80D9DD2E80BB3062B6D577A4A3B6201027B92BBB1D746BF650B766007F35B4ED575CCA11F08A942417639DE2A43BC006857F69F70CEB2B4AEBCDB914DF48C554B81CDF64BDA69090B137A649BE56C409CC464945896C0937C087B8811B465CBEAD5B3969448D4CCEC5F2641522ECD1A34FD55B3B0672B0F28524F109755583164DC8358FFA13DE28824FB7395E8F5BB1912DD79F5CA986E2EB347D23B5CF1D7C2CC3A57D9E62D02674B7E58D559B260248A6D993D2B0D9F246D3F2CB3A53E067DC0DD58592A3586AC0AA4F369CCDB6DDFFB7779536FA8A01483821F6CC91D0C4EE815A0B7925B9BF3C0F8D5CB1222B67CABF5C0A17CEE936194EAA4C63947A4D060158C735819D5BC18E632031A350F384848B46DED7C546498F8D16817B4E9F2FBE000115B0EC56063BE1DC1432C5A6652CC8B134AA0C07026E7721D7A397A26B7852F649B51F4C36C0F1EBDEC7B5C1B164B9181EBA1782B549B635FD2316F726BFA4C9F4760B1E44E66C4C2CC150B9A47545EE9ABD621041476D54D36433A20C1DAD2F815936F65354D681CA59C9229E8A9A30C62315D3EE26232A6D5E721B6737A6F6E4EE443FA50C12AF9151366471DBB346809BD9B314911DC698DC02650368D301BE3BFD51D11ACBA0D629650CECBB0670C476833A386532E240165A71ACE9D9F75E2320784B78BD04D5121847745EDCF24DAF4FDD5F3124DFB449CA8E1FA1B2EF71D96BC8AD531F1353E36C5D44E62B0AA579125FD84AD1CAEBCECC6B8C10E7426F5C2DA069816B5F0F272730FC10AD80B4569F07E3224B9F79D44919B32E3B7B14696DF166E0614480F68224E94B9F35E87F9AC88BFCABDD4E9480CAC5EB55914C117B9B4595FF4E1E2B038F009A33FA9F0F0509C0878D9004B387662F7F6F838683'
			context:   '1C2CCC0BD9831A88AFE58FE30958744EC50BF5695EC031714DAD5A8DF39C85C3DE8F6272300F4F54A5C2B4AE0D0C787A4CA3D60FD5F66B7F9FFC1A28D8C04A63949CEF82D2C0F19B1ACA60C940D06D67D6324D3EFF1A5FCE12353222AB691F068CF47F7B744EAC99E2D62935C47DB5D11EC592F7C6D658141863D07F5AD47244FF2547F5A28C2D682A1415572E7731E3B48CF6'
			hashalg:   'none'
			signature: '409C95E50992D0075878199DF7ACC38B1188D22EEE74F22125002DECC37EB669B58A10EBBD1C3F82B147C7A82219C157105CF2E152DD9583861E1E76FFC1C8D4D92FBAD0052017355E87F4BB33705A3E1B8E8A20802B482D265AA5C4A951A7F7233409F428ABBFAEB8DAEF864170BFCD1CDD8824D3060552065889A5DF490B74523BA0A3EFD0F11F6738944B087738F639FEBAACF39A43E5873E8B7F79C1228095E179C934AB586752C94E63DA65C77507FA6964D16837532D2CBE2940116A4BAEE46AA1FF0781443A2289CBFA0736D49500959002DC798B21D88F43ADBA59C956468B055FB980EF0063B0CD944C996A4EF3A9483F0A707D50070660237BD6D4EF8DB7D15838306E6C914DDD02F0711AB295BBFAA6A8F056A3C7800AD2934E5AB0820E728058D51DDF7002E3E870D7317F7E0454D5750B525D8CF1C263430A8C82CB4475DEFEC93CCF8DEFEEC466E055B4BCF5E2AA0841C601B3D79DA94C7CC724B607723F7A0D6F925CEB7B285BC0F77D026E3337050E90F65C7659E1CDED1CCF7AAD4C45656CC71913487441F10C57C0AB29F1A208EF01FECCAD1C5E5E4E429B3DEE07C2CB71D9734CDA593F662C929F279025DC906B28CB01AD7662E5D5F8A1BE628BFB41961DAC1D93942C87718F247E41B90A59D4A480AC60D367D89F355024D7929048AA8A782E59CBEBF022CF8F6AC2B99AC24EF631F7A3CF7662D34206E5B7B35EDBED1ED9F98EA36C8EC46907FA52E7F5F4C17D8C73E7B9F615D7201C6125E3A1CEE959B0DC52DD729351063E27675C04456A978CB8512CFF0AA1779F5176C4AED38C0A90BFD442A6AE7D3FBA7563FED9D92B46CB541F69FCB0FA6218C56049857650491F07F8498FF567CA22359108F012E260FBAFAB29A31F7C7015C05F1DEE7B47E36C8A3E8E816AC9D46A4731A46E664FD441419BA7432A28C370C83E6BB54FE30979FCA143CA3AB3673890EC101A979E2E0D2CB0AE43A7794D537A9951ECB9A8B5B7ADC918DF8865ADBE4C1CE24DAEC8B04DD1BF8B5C2823854D07D8DAEFBE60E7962D79473B71802D2EA15AC03735B40ADC8A954E791C6520E84075C3ED7B19C5B456AEF025381449D2448B360FDE9F5AB237B87BB758B85F1B470344CCFF0BCE23DC4FD95882C7EBA2694C5355E233BCE27C599DB4F9C821D7658426C2AE6EB38AEFAD52B0CFE1842F36155392A1EC0601B6E4C53D6BFF2369D621633EE6B41446967D473C6CA368D75F1A45D63843CA47D670BB8D9EA2B28732FF979A842643A08BF6E51C0709DACBB617C112167056E2AB2D45FC9CC4D83BF12CB0024437CA98A03C5651253CAFBCC2932FAA160974BD2926AF7F8A5659DC9B9950C77E28A3EE020E1BE610B6BC2AE88F7B7DC5331DB9F7577275D55FBE14702CDAA3AAE920A3E3A45766E8FC6746534D7AB7039F7EE32869127A1371FFD9908A592CE2527E7F2F238AF20C4EDBFC8E0F54B12015D9BFCD4B89A0CA69964E828CE54B93F1A2DFC2D1296DDC3233CB836B08C39B431313ABBF3AA0F7962F492C95C164C4889A35CED0D3FDAE6F3B6876F4C1A069C6C8FEAC8156AE26634ED4297753AEE5D254D2589EB0132FB1EA47149B7B696777E5D41714E2F570EAC2F4868E7E783546852985EA4079DB4AB7C884A23819A78314522868F7C078D2A00A88440F14BB917D94AF7116E92E77E80D927E49615B107F31FAEAECD35E9398232F992E61BC0B23F5882B434C65F038ED1B3BD7D5567908148E477BDAC0564D1B6EB2AA8430924A1F207DE0998B4140579D0D1D9D6CC3BBE071C215AF50E7B3372BA679717F1CB4CD93BB521E851A2674B47FA63A4FFA8534A938214C59C530F902CA78EA105C1C56D329E4ACEA8C08499840C68F6A167481CC072340E6B6844F757102F65579E5A2AA22606F18DB616B26CDCC002B00979D17A4B27AE5614F1D4865C35FA4ABBB42FF3CF19ECD97A3990D55DB588E0CEBF7C4119138465E7BE64D8E8306CD240D8A3DDA805152FC65BCED894B5082653FDDFE7ED79B84BD865EBD341D8B14F2C75BFB11B56BF95657E5548AA2EFCA238D7D9D9C468A9A1B76365060D22FB1C98169CE181C900334C2398EA34C31152C659565634847D90FD62BC191811342D71E22314E4B94BC4F48D767C8C54A3D68C3CF9A09566D9568EB64B906DE01FE2E5FE996DDF0FFFB874FDA7BB771671A446AF9C08736BFD2BB1A7F168FEEE46D422A72B5C62F95B01FFB24BD96039C72FA3EBF4A5EF56EE68BCD4516E3C08898725F51BBB8A7B9B083FBE47E3816A50ED5DD292278BC69E8AC82111ED3FAAB24F54F9261645A07352D8DD8F33BD20859961F076BDCF143D1360C410C59BA1AF4363F72B664D911321CD3F1EBAEC4FEBF3AF2D85327B869C522C2195B05398CB12E96A32DE741249C7B96A2A6C3D6E417A12A8F6D21E104A40910DBBF4960C314A0218EE1323D83DBF68805405D5A69AB4E610EAA0FD4A624AA963314DE608BBA1DF1EE1CF0F070192BA607BBEC877434FA817EC2FF6BB3E6A54953B7505DFE26D9C9E47078FE2304792CBA4696C602C86595627D76BB9988011B70231FDB6AC64337DBF6269C57F285F36F314E476B3149C9B43C0BB3293A8CAAD54AD84AD1A9FB5FD4167E17FBA4B92B1CE9B0D0E27342142118375A0EDC8C90E2AE4500305045C8C3CEA685F17E2ADE2A997A49C2111211272C125F5E1BDB279A7EE355281C813A54B7D662DF62AE72600E2E80928E94F0856340A3C229622FF3B25E1FD2E8578411A8812928B07C2654B409438492EFC61AD38BBFA4631A4E6C8BA6CDB7958267F2977D98BB4BE4C9496B0AF0D688D989F8BEDA0012D7B19F4309AF99849F31269F07602123CF73C77D7B3ACBCB5CE5B3B80E439F25104854CB7222996EB72584E2DA673EF1F3668E82E3DEF0B1D40F8F5D8D3A97BF1538CF19B9268B679E16BFF5C24A957D898D7B84D6D2DA4A11EAB71860EED334570DE3F2818A2C0AAE180014EEEC02E60A9D5C1FC707C6B266D8DA7EABAB9C3EEDF29653DBAE8875AF182C3DDE53D9E0A6BBA09CB023F8E4987EC7B57861BEABEFAA848EBB511FD2FC8D32B4FC5B6BD77DEE1C6A4A9F2BAFF1B5F8B0E87C5B62F712DC9B58C78A8E46DE849E9822DF86B944F705E327A03B91CDBBD759B9B95AD76F90D03E4E2FC155C25C60A87F0838C1A3E54DB09BF5541F722F45737E46334D016B12EECA232127BE99D18EA5D596C26584C4442110DFD2610645E5591CF19161311783220DD8036D916C5EC6303C063E8D29EE3A63851DDC13D00648E32A14DB9137087B9ABD615DEC20EA1975FB9514B2999F21BEBEEB889C2C1CB9694C98FED685EA0164690CFD09C02AABFE1F11BDE56780509AE622A281BAEB64F81DD78553EB51418D21A6CFE805A02B6DAE53BB4CC2AC775837AF92D617173EDF8440A103BDA0AA6EA7DD3D2E5714267529D700B7A74FC0350F5D4FC6C4A6286E5D8E2B999E524AACF519B24E7446385EF645BC7056DDBB0EC071BF5196B944DF7C681AAD337E63A5D1AED7AD59FE329155EEA5E81BECD135DE46B04281CB6E2276437F814A5673DF73EA5909174E63B249D20DC8E43A4B312608BD42DA8472492EA0460A259EF753D479C789A4DA6CD95F609667D9DC48B22DC19BCB2523B422C739CDA1B57372267A0BF78BA7554A116681E1E899EEEF4A08B9FFEB30AFEA5C8355EDE8C3673A6D3B0B5C685B0F201755DDC2E34C2D103BD3C3EAB2C178C5529E45D23B2C8EE990B366C3BE6F5800644CCD3CADC391A44672A1EA7CFFEA1672321FA81518F9508FB0C630026341976A942FB49044118D5630317E32F0F647F14532AFE33F499AAF44F144930E7F618A0DD9C94382D4D6BE999B7481172FDA5A07E43824E2A6E91E30A7FF26347E34EF58AAF77F9EA88B0FC63C3C732C505534A0735E0DEBB9B0F6C1E028FB0EC0EF8478AFF58490E51BA9CFF934FD6D79CA6C40FB768A6F0B8C70F9BC19D18BE96C4C8E451BB9E858970243242D15961F6B1293CE81CC9532625E7026D4E0F1FB0F66F0938EC94204F0E3E43B3502F35B5A90601F133C2517698509E62E8381D3166C48785EFCEEB0A5A7672F91CF31DFEBAF928AEAF13460B8D5C847A399CEB1B9D805BD7270983AFF19759CFE2C2FBE78511ADFE8DD6291D07F66C0F2C81AA59D509C94CF1BE40EA2C0AF7301BA3D0B8934A19F47265F8CB550623756E60E90E3A6880BB2909F1E5734EDD88791BF6DADF42029438CE0CA1579E22914EC59D9516F1D46A9EFC791BA2027BDDF39446ABFE60B7FAAD6D67F8F31D87E5F2CA6F9B89B42D11307C69E89C36BB4090915D07F44C0F8409026D86BAE156E3BD536ABCDD3AFA4A8C85F4E06FF78FE0631B945C52036A325510E9BD1667478B33A5AD94C99881CD793723B83557286986DA0EE7DCE46C84127E60B0ABF7B8976099D3F4F6AAFD7532FEA52AF8BADACDEDD367175FD8102F5E52BD8B0CA521721A22B0EF4401C2454DF4E361CC736D3230307D5634B0BFCF51BFF9ECF769D5ADB772D5B8E91F6EF44DB72291AA5E8F8C884AE2B50DFB5C14840344E1EA3A0961C1EF20DC274BC8140B22E13B4E02D7B690856ABFABEBD992E0DF8261D5489FB81DD3FB2DA64458D41B65025E14E468204E028E38F2ABA3EA55E905CD5637EBEDEC2DAE224277C6614324F598B1602C025AB46A62C0BF157B329533115A6098B208916CDE8FDF52C23F297B030FAAF668D2DE50061282A2AC1CB1D34911F80766EADD77157D7D7D2BBB18BE4AE9D8A97A80AFDB10D7B41D40B1453D65843E2BEC623B77D6B8311A2BBBC0F57BCBC6B1955993508BC2BAC214403043EF641B7E3004633CBB9391B5E623615D7F6F89693872BC8A94FA72A05BF4B836E8377F9E04FBB347DCF7AB11243324AE1DBA42A0551429E944496ABC4718ABC2840878EE5EE9EFDDF07B20AF29219F7BCF020FCFE02EDB05E6F97F4BC683B238D28DCAE65CE3CF2AA0895FD3FAAEDC242CD66759449630C73BC104546C248A735EAC833CEC4D5E2D05C89D2D4E40621575877FD47CA1A0274A1B6CD7C4E0AD783B1C5DCC821A7D7D33F47F722345C79924A30BA0A5E85D265320CEF130F3A5237EAF97F57D55C4D57D48555FD654884F3F67F4FEF7D4720148921DF409C27B6A4B18CF9C3FF4A9FC7B4B30F3D7A44EB6615FC4C54393827623C96A62C1BF70990A535FDB9D22D3C6336FBB34B0549312847D5CBB5D4A251088026E169A5B7541190016CB9D454B0EE9FDCA89DFA99C3C1112FC7A48C720A1A4EF767D1492FC335D0D1117DAA3E9783964EC3AF9D363DAFFFFE07ABE1276AF528148955DEB3F6FCB7C685971E4335AACD74015819FFCD55104493806C3E4CDCC7B55DB6B187EDE39C638BAA965F25C22010888A9F6CE4DC81EA17735013DCB5E00B753A977D910125BD5DD0DEC878C894FBDCFC344B51033B00B24D6E43C42AEB910F9377AEA0E04C35D83E89221646110365C44EA35855B1825AB6BBBB3FC648BA1AE5EE2FB1BD527A128B21E9AC8D1298EF6C341A0A0C2B6290B00B9FAFB43D6CA5BB9B1359CC4B6FA532518DF5C76BE2AC003ECEA157CE987071ADB74B1A61DC0D6DB7E71ED82295336583642156407C51D7721FBDB3FA0B4B0ACCBFA57D94D76545AA787C2DD1F9F82D7DFD0044368B2B092A5B855BA6DA394D0AA84680DE95A3D8C332C1BD5C3D2E011DB1638DBF2AB26E0FAE9FA49F7C72C2E8B384B7F7E784E2D2CC9BF15ED81D7D19F5BE2B7FC23A11E69146BC155D6046E63A991A3B2E65C889BF4B4FDBFF125C2C9EB97B509E1AFC4FA3A6EAB399B89518FE08A7A262BBC04EF1920342F29F799D42DC292673F051783983BBFCAAE66B7677611BD86A7158AEC7872EA13DCB566995DA591DCD956155D3B85FC596CDF3E3E06106C734B915FC5C51CA83B9378183596703852B150E037221A25DC1795D0AC77AC6D5D0684C6D292E1F0B887F24871D22430D8AB4D9C6CA34D635A13FD0F226C5304AF6FFB560CC3D3EDC51D692EE6EC907F7559C968A990EFA80966B4613B02902709DC53796F4B07EE0A343620A5011DA423D22B195D8BF75D445BE31F8AD0DA51F0DF461758855C5838C921403EE43D366324EA1F65FCB6916D568192042E8F6AD9589B57E267E5840B2ACAA2D3092773F98968AD9602C85C4D41C1DB32E842F4DBF80F2C5ED5013F5077CCCFC55AC0434174091FA62DDEE627CC488720907AE0EA31CF0252D49DCA4EE66401255250A53839631697E5E8017E349D24001D4EBBA9C1D75A9E9254E8131F02C0D0010AAACAD389EAD31E50B290E1313334784C0E28EF90D19651EB4DAF75215E013D6D569366AB211D738A5F599D240AEAD9FFDD014418CBD1C8C6DEE07030832C134D26E5EF960CCA789CDD4BC29C6F7ABF50C03520CAA39CA07D823CC7E4FF67F6DC98E18596D273434DCA47354BD0A9617C66D360B018757915472F76A87CE8A4979BA9B04864DB95471F457A3ECF23B9A8BB889E038B59A4401FA5FED0DB83A0A285161BF78B503E9D9651B8E41FB39116FB6FE2A5402EE9A8A1C145B5B48B4BBE91F546F3389B0BBDD4F83ECEA4F00A3EF03B029AD896ADAE1F377A2ACB8B085AA91EEBE4F6A66E2E528940B4DE228B21FDDD655399BF0F2959B19DDF9DC0BE17E0A812F3EFAE77CA73F624F42DE87F8D255AA90B7354E51181C6970ADD37D5220386CC7728CDFA3BDEBA13710B9064F1D804E22DAFCD69C5E58B20518F92A69441DD5DADD67BD5507528B5E792433DBAD7377676BA15CE13C454392FF34EDFC06648494A35EFBFA89B67CAFA06143D4E4069B03FAAEA4A6F9C85555689EF2774455183D3CF4D7B3EAB269873895DC37F4E9C054540C4DA64975D0FF7A68F37011EBBF61D4922154F2333E833B90FFFF85338DE45D2550FB84BF86FF47054538A921B123D913DE8FE30F7BA8D307F195E3E3C5FD4BC49878CF22807AE18FD4E3E05B5B8CBF6EFAFE31F3CFF1CE9978C09D99124DDA864A6877E5DBA71FECFBDC07A639C97CA6ACF3801D268F2F26926CE21BE1A9D10F744B4797AF8B6A0CB5E8758C84F9D65929EC1B6E6B6B09082AC5CCA02DCD7B088C4FB3892D083BFF44EF090CE09D9259231AF74007C72A856D80B6A51BD5973BDC3EBFAE2CB86BF6E7AB9578C82F69AF50062ED8FC8BDCFB8FD0B82555838D34C273ED78C121A0600EC860A7816FCE9DBCEA227730CAF84AC9BF7BBD568E46CAEC22810CF456B797FBE2DF3B25C73BA81498587BB18FBB5E1582E93B2308C6C0C34745AD07DF4AADDCBAFA6F58836D82A07159011B82F88DD9B36A60366907F941885B30EE9C09FD31677AAC82D81A59A1D9D0BC57105D5D4E45ECB19E3E70464F791F76D4EF2FE86D176D3BEDC7F33701689525802A129FD92BD0156CDC8539D76F1B3724B8B9350DFC6587DCE46096868A1C1C60EB4C1F89CBB05AD0D4EBDE9B3DD9B1D87F670472896B75064C695E4B5A66F6E5D4C1EB217800816C8D1319B3CAE54920A618BA6DA437A5019B53C1D4A5D57C76D6ED3AECCE3B0A1C893071B5B97FB619BC4029846B8923632A49EA353E70B9AD7F1E44FC89FBB60245837C9405530F398401CA973EF5312B1FB940E06C1CFA7BD5C8FE06C1991E9955DA1406BA4E0A11ABC3D65EB65A24246A30474F97FD164ECFE963D4B705913A8396FE1C08AB46EFD6CE1C7A57C228111F8B18FF23320E7EE221B17C35B3E12226D756F0FE7E831B84D8245FB731FA9188CBFC86643D6590970918F049BF5994C0B2742C7FA8148B013BDF95448019F67C684D9E31AE501DFFBFFB7CAB7273D4A00C1D081B07589A6776DC2622E3F766EF221A536B971D8966F3BDC997B48596865DA12911F00FA7747F9D234EDC407DECE393BC2BC8D1B5FF35B38BFF77C3A5B260CDFF0205FF00A31219EC4BD2C9D162E62CF1EBF3CAE66F73F5171DB1FC0DE595ACB1CA1FCF345936FB9B697F05DF6B1F725229D099C177A2215682E68CAA4EA89BABF101E6830A225A1D56977A8A2564E1C16C791B71A46203DEFA9E28BDFFD1B7893F2DD06C4FFBA6869158F721DD7ABF01B450B253F02E53161F84A67846AD505DC98C70718B65097CB71D1D5F6E6B5BB48EDF4807DC4017089636F0A0AA3667BEEC9B9DD9B063D275DE7985E1F9316967D8AF60A0F2EA438944DE2DCEF4E250F28F250D6FF6B334B2D454BCE028EF9AD02F95E78A4326CEB54BB50B2CEC8017EC4820F1681372180D0D5B491C93C2FABDE031E53ACCABAE3F7C9605E0EC302AA6A456F7D2486F48089E0A2A9521EECCA16BA0B119BBC24D3BA64453E35AC58791F289C20B5DE71ADDC3EC81AC45E4C9CFE2C5CF2963CBFAE540672E81B0C8655CCBEDDC584AD029914C49BAB659E8E1337DF8E3BC73059BFBF38F9F7F20D04BB3B0B79134265C34D96EE3214FDAE89E4E3FE427BFCA7CE4DAF5E63DED092E897579AED5F8DD823CE44A5334723178BEADE48820EC7C01CCC8A6D28D9C4ECB0AA75E54D022EBC7D4B6402284D877F830E1C2F361800B791337E53171C16A50D061DDB933E8F96F971698AB6F3CD85D359FBC8AE494AA4C1429623BBBAF552CB5EC8778B95B7E55F34885D2669F823E36718B287DCECB582CBF34016D3013DD247D635F6A26ACE55D448BBC89377E74FDF8AD8AA8EAA87024A55A1434DB49656FB97087BEF7B485121BE354039990F308F9DA6E0995A445C847C3C85F8F0BC48BCFC7F66A960C74AA6CB55E5BFE8EDE100CE8D79F5DF95AB9D082DD93F81DF2963E7EA7D1D439039E11471C8C696D5F74EA13DCF9E0F05636C4145B3EF004F19F9C7854D2466D0B50F6C4794ECBF9CD9109E874936368E4566935CC845B8246189976FD14E080EF4ED7C3C8ED9AABEDAC6DD62BDB7869C0727A5B99D4B25FE1034FEAF9DBE395B303C66679CE13ED52ED254ACD1832A779B3A6A33B05E064B931BB34D3123277C512D795CEB280EDAA53094CDA895E0D7206049538454376F799C676A52FB08293ECA2760496BFFB8EFE3120B76D6D1938270BC224D3FA2B3754EDA7501E1BF71ABE3F6BEB0E9E0B94D1D09208E31BECBEE532C95439075C81748257E029CD3BA2AA18AE89E4AF7357A96FFC0311CCF64A868B7D25D82940A32F7EF6E882A7B0F6C486987FBB672D9A317CD3E9B5F6C1DBB4ECAD223C2CD51DAF054FA65B3C1B907CBCE2CBC3B30AE4776ED98152609E3673E7E1231AA8F4B199F4D42676A1B6FD9FC44177C4887820A6C0AAB6272E9D4720E39D8F7945E2E7FEC5137EA8C3379309580E4BF97C810176678640297532AE7F6289FCBF8203FE3826D8335D40D17A1A3D53747BA21D0CBA617D5DE739C67CE0A618BC9211C42C5F6AE1EB049C4CEE07BF624AD8F6494CE495CC97A7E5A906294A243D39D5C9383632142A3E9CC2AFBC337C13F207F5AC528647CA45916BE93781A16DDDB4E8F14CA57997492EBA2FCFA45FFD2F874C90F2F667FCB1C04CDB093869534FC0A8B5DEEEC16CF03590E789C270E7514355CBB081F823F15DDAACF8D352E0B0FD1092D67B9D4A9F99DE1366737B53E4F477C77EF00F1769115AE25D85951C33283E40D07D18D154B31553B9977E4CE0F848A010420E6F60B3E8BAD3DF1140A232C9F6CFADE4C017A741C738A7E82A9882D556E46C1A7B5DAA287C590EB40EE53E126D7F55AD9C441B8C8B50DF876D37941768E17B81C00840ADEB0A16147C8327F1606A7E2804361F61D45E6CBBC04C7126FADC05842B4DA7CCD4C9D6DB0AFC4EF564B32761248D82F8547C67B895D325AC8BBA1D6F4A0DE6CBDFBEF4C96EFA6D474B545376D94F92DC366EBD3FCDC016865E83F0899137E6B41449D113D3E72BAE5B09C7BD0026A1C9FE4E3F58B35008D6A95896AB9036E79D51FFD3D7BDD2ACD29778CC8DFD52E7C1163C425EB648DBD32F0EEC15E79063D77A476696309464E1F43AAA5A13B3CC67542AC8A729E9520B5146AB1A0929C8FC94760E00BAA48D7ED6EDD5C1E684CBDE3A58C8681AFDB755524B0B79980F20E342BB3D4CEF638B5D3BA47D543BD85475C5C2E8BCCC21E16B7BF96C47265460F9EB67E49CF1E76CF6B329D3408F568E93E52DA1AF2538DF5E431E044BD38BE276DEE8494D1828A89D6271EA76449BB53C74E17645BFE41A53426389C202FBDA7EB8BA7D6BC32D0528F14CE611E12BE32C0BEE52E6447E5E8303E2EA352E9FEF00913E123921FF516261BDC62C490BE377B60EDEA8C12254235CA2791139EC1CB63C9E5D23DA2E87344063918FEFF74B9CB3F98A2DF689D927C472F8C57C2E80A8CC6895C6A8D535A6011A67A45156AC1A9E06C8316A933FC9D0EB0605386D1240BD386456166FFE8BEDCF835E2C1F6B638D1E5B6ED75BAFD3DB79D598EE102F135A0FC7E4AE0DBED17B2EA5C15A0D42C97B7F35FFA7ECC8EEC47C06BBA6EB127D1C6AF7387DC84C45EA2384B6C1A1C79F3AD48BFB92D807AB669CE7C5B183B1F59303DA27DE88055410A0061BD42E0D2AE943E314D945A53BDCD3BA9CEC4D1C767EE500391B93516CBFD517751735E1B4704F0799880F996D1249CF194BC1E4CA2BEF637D39D1671BA0E620F30026B8E3B7F0021E8254BC80C950F1FD53924D3288BB526C7513303DC73AD341F0A85EA0EEF238E35598F27E07920AEE001848AB3329A25C79A5DFEAC647CBB4D557775418C94AC8EBCAEBD960AA44F7C5823F8A72F0084A5C0D485B9D71EFE12E51ADE909D2462E23CD5824CFE6D3ECB95168ED1FF7DBE0FEA860190F606F3C6AC338A188670C343E1F34CEDACFF4D273EAC3A9D72477A2473B34336904C14EEAF1BA384F4FE15570ACF5F97562C713F0580C0188A4830EE48F29875B77CD7A4651AB364E35967EE7FC4EADCBF3DC6D8959B73ABC92A24C2AD648528B0AD742E71689D8F9E63634A2821CCEFC681AA973DA9561D855FFCAAF92E3B8B0A492669EFCC61968093B6D0DE83691B9760863DACA5EE715417D818C3B88D80A650D90AB2D77FD7C2D92DF263F2EF92ED25A241DC4D7C09E78094F08D61183C71436CB259AD309989F123E174E6F6EACF408AA3817A3D2A0A44CDAC06096B264E629E133CDB387E4E7C4C150322EF40E574631EB40560D08C925E0020E9D45118BFCEAA80E61FA11036BA3CE6BB3C86802483285BFFEE094F5D900591256871F44A6EF2B041168A6D292E84F0CCFE4626B23B9F99C17CF8559393F06D536A2D0DAA3E4FEC1B98B965A63A6430A48191ADA59877118A22FEF8C057137203116987C314DAEAC765B5409123827CBDA8C3AD9F78A4B34DA6461EC4D502299D2CBA2DA230458F05F6F421B1C6F31508798E80EA40F6496B7C323F7711D0D103FCB280128DFBCCE149AD4D7BD43FE4E442AA4CE899B639BB72B8D6A93BBA6C4A5A7B07E3E82D25CEF24FBB63B72212D912D3A46208CD5FAE87A6159C49AF915651CFEDDFF075D5549132112C01DB65F917D2D9DC32CD9E2E9864AC50B2BE82F6B32CD774513B73E628EAA59B54F747A5D21F6AD4671AB2BF6F5E1640D5ED6517306984706CA2572BF0082904AF4C8D73BEBFF6BE1CCBC4A3DE0A6920B786D5426D8A69B2DE1BAEAB8967A9DC7D19B10A3280C3DF319CC7B746A96E7DCF9D014858C728077237620B3AAE9DD2629121BD8D3D13B20C84797399C3FA438C78A90C4A80BBD8ACB8A7629593EA5D081974C80AFA81C3E66849145BC3D2765D8DD1FFE14628E1020139C5849686F7AD566CACD77EAD0A69B164174E81546998FCAE3A8F17E28866AB33803BA2E22957D8C3D092A271CAC3526D731501DF0932B91FB915AF1D7D8AC3AA9A0E879719696EC5F334537B137A860ADA0CDA5C4C315B7980D38674071659C2603E12B20D181568D290387BAA91E4F8D14FFF347F836095E9C379BFB97D1E90F6928D8D9B1872308049C6C131F322D6D9EB96D3D2202FEFE10011FC86ECDD3C24FD3129BD50BD7B1510F91FB400EC7D87D1A4D674F681F2908C5679E186C76164CD87DB520BD42E6F8F02505DD0ACD9957CC22F13DD83B1CEDDF2F55B5BA2035D96AA0628A6188B427ADEF559005BA525A9DDB7A4E0C3154E659C1B8963EADCA96621167B4BD18930FE9DCF0B3A0483516F20EB17BF6249773B2CE1A9ABD02385EBEB2E537E8DB37715AADE92FCBC510FA8C0A1A15C72FAAFA493E704362FC6F63B08AB3E68D5CB9A06BB8D1658AEED9801A47DE9239A0824D235CE007AE9D4047C037B9A9F28F99539477A4D96CE5B9744AC81F81F01E87BDB7C99A1B396DA20932CC5FC0E3F402D371E9CDE3239BA60DCB09BEE489D0E307B14A136B2601A6BCEFEFF84E88CE6FABA95FE525BED13B4217C30645CF15BB74C5125256A4A90DE5473DBDB375111BAD116B152F3A6F3A47FA0C53EC88B168CCB59815F591D873DA6D81BE314ECBAAC2A7C7F295CCE9A9B2D4B1E8B27BE122264DCBF6FE467D825AE39F18959150138CA31DB4E002874490CE2AD8034A481A17C925C1F5148547051FDF46BE0CA2DF1C217B7BA22216348A6125570B01BEB602ABA2223D7A17DC72306FC285D1D196A4DD64B90D776F94B83DE7E8EFF76153164085D804E86D785D8C95A79221436C98EF6E246566754B0900F5EC0FB218ED210BFAAE94B7E4B8C3C1A3ED7CF6A6A38ADB08476C43494F752C2B820DBE9BAF6A098401972E02808D2B5F38628BA1B938435C6734560588DEDE49C56174C22642C2DB29F9CC753E1387F1E5CA6B1270E9BE3BF5115A41492B3248649E877B93CDAC58C986418A471D72012854769B549AD1D106CAD8C22C88E424706F6F8B654EE1D6C524FC9FCE9A9E751937CB1340E70E56B170D1D65C128CFA7E9AAFD89BEEA3B33206AB59218D4A103351F4F9B892FA37AE7C188E3D69FC5CAE6A3E321CCA522908BB3ECF347939E3CBC32D2126C7E4825E392CBEB98A1A3097AEEC8A4C4168E27D8BFD3F5F7E20DCEA77C28FF01676DB926914F86A5BF1EAB0F2072490DE6234B5C706FAE2B863DA22E3EAB61AC84F2704B0AC9BA47BE38B629AC1C5E857E92BAC5D4877362634EAC6F86FE839B8E7B8646501712B925085756AB47984BCDB9DECB637832EF106281319CA8E0567B427B3E6DE9A6A2D6A00C999364574921B172530CDE18515C0043C51AACA133413F6A9112348C551427D3BBDC2A546EA744AA056A3C059404811C6491A3CFAB42F029AB15E061A9AD56865E34C287244F559D111AD2349B963D46C86F6EB9391F58C48C17039014684B701ABF6AE358F759630524B38AB6316FCF90273F97FD9C936D77008687FFC9DB0865BDDF3E952ECE40186DE27E3392139A684610FFC91277AD2BFBC2EDB644836B75499EB8F176F875A6CA1CE733315FB2F70171A21F6F43BC735B8BD06C29B30C6CC5D4A791AEA3C1246CC0618131A07868916199C783BF9B85EDC6F44D9EB101D274AAA391176835BEDE8D1C493F85D07D27C8CDB37FD951825978190BF03D343B354E6F7CD48171778DD167496A185FDBC654F315629B43347F5A9D3450A38D16B1D22B91E30FF3B77FB1602111F140DBE64C0B34B64D6AACE20D1B40B938EE1EF12968C59A22EEE62FDFCD36F99497DD0A6A3214B7DAA23902D5EE3389C3228577F9D34380B3A9AA4B5354F959FCDD7AF2FA7A23D671987DE8934AAB537B7F79A28E26900B4B4ADADB2CB37A1EAAFC72CB3F124D4E723597597D334F799E8C66ACC47E8059BEFADBD7EC26405A9F98FC3340FA261CB072E4EE15334C1801B7C7654CEDB70A0CB57B1D0EE2E6C9FEB8A0E54C195AE275A5BA438FA12B60E15ADE624667DCC33A5D864354CF61CDE232523E56974A4AEDD11301BA7DF67CF0B87AFB5B695DC90C943EA08C1E75A7861F6DB74482502DDFDA7BC2F66E4AB1BBF1EAA75F39638106A97FFE7928E844FBD81DD2A212D856001B15F06714547101ACEFBDAEA27AE5BBE461B25DAA902D3669F83E4ABBD44C92F047121E9ABCC8F3B340A8DE6346DD1B4F918BD72265720EEF2150DC6EFBF058DA6FBA5653827780A704E513CF03F3B09D935E70CCA4D44A077689BAC59EFDEF8FC28B3FF0D6FDFD68E5A212A13498B091EBF0B2AE5B9926AEFCA7E76260C94E31EDCBCF5F0F6CA846D493A0DDE854CF2E5F1BDA212ACEDFDD3817FE4E47C6EB1675FBF254F096B957031AE90FB9AADA2266B213EFB54A17B6D36717227E40ECB455C18C5DF72175BF5BBD26F0E7FF89D065DD4D5BCDB6DCC0BBE22537326125E2420DA31B1466ADFE49073D33EC4CBAAFF7E907A4EDF8B777D6EE579DE331768EE8844B89A5CF9E2776AEAEAC8AB3986735B697C54D2363E74B6528D3373AB0720DB55B315B73B8AF86A7EB486D331132E18A224A1341383275FAC663F74BF0F5A6C581E63EB60832CDB0AEB99C87C98709178DFAD7F9A08A0B699E47D5A14A8A344032C59F8412F724BD53A5300D73F37A4878547AF8D1E31A1CF399DAD124926C7887B6E5B0DBA463398D7AA0627856ED4F75FEF9CC27546289E769F315B8A47410D52FB0E4ABC89DD4D46CAF61E7F4B060940ED87787371A016AF9DE6396AEB6B0E6017B9F8F10FAE7F7C3A012206BE75D6F08D5E6B5CCBD111830EECE17AB1E297C41F820797A413B73BF309E78082880DF6FCBCAB9AB08E2362BDAB74420322EFB4F595A5FE95710E95EE1973606FFC36B17A2A21E5FDC443323A1D9F72001F86523A440B82BF4A0A5CA71B91CE9E5A788EF5DF93E988B911D18ED4B8ED5B184F9E09DFF6AF6A95BD8B11C914421AC3AA7FF18A47F548840B19105DA2C337EE94170E1D1A977662A611C3C3464A11A5B0B918DA7F29A13796323D605FD879AE50F843749AF4F92CE07422D60E377788C3A6EF21387F84DAF8C40ABE66FBEED8236115FB6FB7DF27294EE58DD7FBDC1B924DF843FD165FD2F4E6BA9C1F2EF69F354D65BB29A9602CD5AE2897193D77B8BD3E9E64AB355965C2CCDD575A9E7900147EA7693C93D59B13697C6C809953FE648E81AC333989B0850F42CB2837671F8A9C6D98B49E1BD7DF2C241B424894EB8DC51D91CCC259321B7F00956165654A4D5AD3EA560F5D4B1E35B3DF1EFC8C961792BC0351802B1C5032154DBD9FBE3A8FF270D43B663D8E48D6CCB5C41E71AC828BD7ECDDA0090FC1C663A75EF38030F1B6C7FD15BBD330F37088E61208D03334B74AFC7EB17D50EE6EA35003761BA4D7C6EED2C74FE32CF0CF91DCD8771FE4AAC3852A41656542715303BBDD2F9501F8FEF0946F8C8E352B8DA664CB8831344A3C8EFB4B105C48E5423D53151B5BCBA390EC9E28DF3F8FFCC74FC20A5FDBEF58D03A72003143A944CC9AFCAB938E8A6D755F9296ED2A93C97FE3BE0D490A3F1453B953D9B36E95F7B7999E1BA3D93AB27600700A339B3FDED48F2180676A7EC75121D39FE87161FA28DE2C27E1B5948FAED3E6BD17AA9DCEF29B2BBE63B4DB3B9E9794B5F6BD53C5562AB12879823820BF9A4741757832675234117AF7386A6DECC17949A2733FDE7FFF3C6441EAFFDBFC88409A19EBD95BB038F222E379CE9EA54C659FEBCFEB18B95423075C726389D953A224C0B2072470F6AA9926D3ED5A0B755EFF9FD236923B7ABD191A0443D8471BD43010E328DD8510D66EAD7D9261BAE47ECBF53C9EB668520038F66A8F327E28466E2EA6D4545E8BFA9157DC15FF6DB39B14E2193CE2F475C026F32743704C1D095497B071522A2EF3E72B2700677B505E48255C450C9FC25DE6FD1D706D8D54CCF19DB6F7447D8623C6FA01B2763572702093671EC0815B3A41FBB6689908DDDE9144B01AD22FC6B1DF316E76848DE9E6BE912E69272494243DF924B63513600D5AFFD3B1F07731AE5FA3692BB0F17720DFC60D54329F362D4E0B58051CB757522757013E4FBFF3F8812E6F4277261E6BEEC836A3035EB21D154974659ECB5E467E09A331ED4DA4F7A09D5E411A984B909D6B39D2BA1CDCACA7EEC3F3F7388B8A3DA655D4E8AB8972E1F5A3930AC7EBCE878FB24ECB496423C2D013BD15528332F5060B7CCD274F1C784DB90A755E92A7AB5B9DDE9B2FA40435412D978C620748EB4943A712D2AD4CD35124B410FA7DF07632F22A7F6E0E8B8FF74E73032AE4A26620B1D441DFCA1D780AF03B2A255739B1F4CF18679522ACBA2CACE50FB4628B04FCBE9A3C7D6B1B11320240E98501340A183FCFB50734F8DFB95070876CEC69409339F56DFAFA42EF6656C5F1FA55FB89AC29723C27DD44E793169AD3B0D916D0C7E850518C8E766AAD632B9A1DCBC47228B6B2E541F890CAD3A90DA5E6BA86064E3D61122A30BC248E3BF064E75E19C97DEF616FD29DB66D9680C9EAEC364B726AC3C84AFE6F66663475B98C427815CE36210B1E346E3A271BB3464522198E226CE6F0364458D3049AC02698D72119FAE0C428AC7DB2E34F3B8294BBEFB2C3DF3AF59D9B42A4B4ABAE1176C40EEDB5B4CB2AFC964071490400D44664D9944179F9C057673D679B533C6F69C44967AB9AB3ED2944C2149B5F7B8A09408385E46199BECFE48E74B2F7854A09532383FE46EB21C0BBE15EBF0BCA55B80C7B250128CA76B0D3FCBD13398C7B43F23F8DF2C27E0882DB822AF3A77B4B2B8708FC6924BD1CB9B4D8454E4BB3E3A7A53F814D20F9805533B1BB5CA126B63699C96DD8A90275F10EFCD87BCEA35845B8E9A7B1A08CB6AE8719AF095E631ED1B4A341BE94581627E2467DC53ED1CD8CA2CC6D5142AA268B17515DE58A6C2F22071B97ADF8A2694F82A219BBCFDABCD34C8B78C29256DEA19175460450B843F2459BCBC6E7849C0231337DA5C62C3DC650EA762239FD8E6C88624434F82EF72CC471686DCCB14DBF063A3F0AB8FA70669B70067A03CE43E27F8CD14FF0EF12CDD26F1260C8AB54357A879C347AE58EAA2E489F52FFEBE93C37C98A72F470D01CC6A93CA2540A27173E86EBFB7FCAE8F69370C307C0BE10197FE7E25F0776681A01ECF3AE7854F54733544710912574821C8BDF8E4D87420A40934F3C8BC411B1965C1B63C2478564A12B123D687D1E8DA3C242827E7B81486A5CD973F0DBDAEC4C9DD8E26FFEC4B114E778D8AFA2719F0A3223EF8CDC282759168A545008C465130235872A38C228DCBCFF650499F780077B3835A7325B1784AAF554E29DA918A722D5A960D380FF898248AE78678B80C0C90E7E248D87394D166F5F577C997D61242B0EF76B181659720FF819E7B9FB6CD8B20A47E2FCA3FCDEB0A50A26CBB5C4DC382FE7154638D2A62477CCCA65C5F33CDCBC9B05C821C0463DD6729FBFBB9D5CC461551B4D0E508180CEF5E44C642853D60C41FEE37ED02683C242B7E2EA0DC6B49A8683C3623367DDB5F179A65916A192B5262A393C0912E9F200CF638E170DCDA99CF4863253AA833737486A7D8D257D3C8418DB25070E4AD1ADD19E1B8A0514D354227C46C5753EA93B84C27F865DC9A6A8C398831796B478EC2E74A89498B516D2D5E3E38161D6A62D5BFDF4D128518FEC54F7B323840A36E004C56915E8E13E38A2AF6AB4002599B45F820A151B69B853993D989E08C15B1F698F158E377151632144F82A47DC125D1671D875A61E6DDBD8DDD7CC347DF144EE57735D8A5D669F3489BA1AA3B0D6FF6AE9550FC1F459A9E159F659EF0140C302B04435102AC96718A0C543EFDCF5A04B526A56543BEF3A1F8C3EFD8430D90A22460201541445A2A02DDF70E12321C986CA19A41720E1323D007AD18F78DD6AE24B43E119DCF53B38497A39437E217B0D6B6CBADF58B9AE45C46DEA630BB9D720DABA4B46C85B864116DD390257BED7450292E84EA5007845429562D001D6B388AB80E21E03E2CE49788AC70535A6ED37AF2033A4B75F49734A776605AA287CF28237AB5F8BEF1F6FB37F0DE6B562F4A6A43C0C8778224451796C0817FE94E02C0860ABC48E6790F8C61A617FD4401F838C9A478992A2015FBF64E5D1B554EDC10426339F14A9357198AAF754E4284DEDA3A3DE7D0072219F2623705577F0F26C9E54B53380CB7226E2C3152E6BF0DC1420BD50A999FC33ED673EACB17F1EE36213371B5852EBE9A15CE607D946578FC8DCA8E94660BB88ACD518D5A30C253801C6AF4C097930A66E4398831F0C00E453EBB01ED143A4B6FAD37F898FF46114380C2CE6EB24D7EC763648C2AC94D1C37836879F36D8FD00EFA0F69DCA05D6387DF3C0A334082783B24FD958903FB124CB6AF6535C758FAD7FBA63F4A549ECCC2833CA7335A3FBE89B61418B5D912EF4186330C9436090F433B9C4913DDA0E7322B972447882AA292A8DC9AE201D6E15D7281D2631DAC7EB654AF256B42255602E706D83B0A2FF2FB7A1634798853712BF434CE5A9B6BFD830703A1ED66D7ABE4EA11D6DEBF076E33B513BBD6AB28BC0F9A79B488EB8C6594342C713811A4CDF657B791751B7F0F67940179C473B48FF152DAF8776ACA61A1757A1AB713DCCCDC042AF08BC6B7CFFF5F9A3B78C6B0E728E2BB7FD014CC52E47DCE0930BC3CE466B757251B6EC0A00FEA5271C5518DD1AE6FF8301CDF8F6F70F43F709B98251F1A910BA06A2730B9408B32C7BC6570B6CFAB45BC74B5E7384E74EBDAF482D03BB71E0232F8289E8B6B326A8A9C99C459D5F61F9BCF84A8FD637A837E897F46FD26FECC92D0936ACB78DBFFAD6272D904F39CC34023AAD1B99E89C3DE58AB66CC7548B577E3047C6464C09F9C6840F01BB0D041F6EFF1362163805321AF8A6898B31D16A02FA4735AF4D9859E267561EE8F8AADAF3E84D19111A991F6497F9DB92A5A4F684C806CA84A189AC09C7A3681717EA0031C087BC9DF030E09CD364F644021160874E3A7CE377FE38F3557377CB99B6D41310083BD55C1DD2609F0F75EB0B7802161E95C44DABA5D9FD09EF67B0E508B8E06A91CBAB99C6624453A446791993D32B9FC61CDFB5B974BFAAFBBB6DBF16AA75C997B314316F486F5C4CCD8136DAA0EA2A2222931B4BE97EEE8381D03280EB3D8F83143DCC4FAC996908A50043AF00FD6F238222632BA67BEACDDCDFF0B42732AAA81975EC0D98E4354315CF96167760DD105201F588251AE72EDBF06D9CD80F826FD6AA7A6D186B1F5A1798E8E9C29E2C26DD6505A8F1FEC421CCB5E149896CEF6C934A69B9DC2A2A4A90136C7A1AF3CB02FBD31F6C3A70171D3BE3D59E03578847D6EC738E54C10F9DE8459AB666983DD9F4AF2EBE65DBC1B6AE3F88D73D5C3BBEDD597CC22EEFC718A0C25B5DB255257F493847AD4B85E84E44F67F69FA0D9E5E2E54891469DE5FAC047E13BDCBA46D2844DD9ABB408D70BF8668B74BEB7D8A941B56DE571E17EA3D8F6EDC120528933290FDACE50E59D9001DDE1AEEF5F2ECD14BC37F240E0A15BC62890950EC7A3B7E84EF20C7895D428ED601920717CF2D041AD16FA0FA054287B66CD3518DACBEA1AD8A5C35D5C695C26FB48976D997CCF503BB71749CC980C1A02DDC5D0F9A2195D52767FCB2037AD285ED466264A42C1FBC99D50548338993F8923084C60673ABED5FC0FD9B418B5653FEBCFEE723D62C92221F88505EEC013CDD18043059610B779035128727654EC4FC384BF8DD591342F7364B435681F6180C00114BEA0CEC53779ECF12339A2035A3B24AD1D6429F4C0AED1D6DF61B5A89409E73EC2DA623CFBC955C976DFC9412D1249BDF4A871FCBDA5557E998FD766C413BA7C1E8A8E909B296A4EACF2CDAD85AACB808E54E0BB66247D0ED8925E06C49E99CD1F61B492F53EAAB52858B0AEA1A8B7BF87F1DCFEE24C9F61E6C573A438AAE8A6B56619A5E4CF7ECBEB7CADA7691C1B202332D764450768716D4B66C8BC83E570CA4A11FD10DB747A98AA1EB98E82FF7819A7ED39F0DC55B779E1A8B932BC580142CA6FF64D08F96CC63B63347DEE7674361674C3943776575A76BA55B8AB44C980417DCFE03F96DFBC95981B539B7E8E0EC4F8883620D87F11F8B1AF6B2F384FB65E84488B28D1D037CDFE6829624D7B8F3372130833C4BED1E32EED378D9D0DF92C33260B95E4A073E9030370167AFF019CF423F7F6E7195FE368FE03CA3F362982BF368693F90131762CD61F949A94499210D44AF32D8A302A993981B601B789A45FA5C76B5251F02907CB7209CE646C1947F6319E0DFBD7AC3996D093023EAC2C71AE61E936FD7751E31A594E0B739A010B7143E86DFBB1E62F0B0500F894D4F8B44994D47B74F8B04947D9E061DAD21C96775D5554EB2A630E0C6604EA82A5E9F5C935C3E807022F28D033EEEE52E570F9CB95B461DD6F63D299368BE940EAFDC7BA888C993639F75ADC2D071FBB99807B6E420C56BC3BF5DBEA3FE3D113A9314DB118DD7BC801EF8087562BB2266332805EBBD6E50A61EB2317D504E27509F2E864A8C1897A94995685D2B01DCD6648FB0259620AB6DBF1F22E3988A6EE5DE4929100653E4B00D641998497D86AD07CE32D434D395AFA535346B2C71A4EB5B9AB1993611356FB80E0EAFB446FD19EEFBE89B0427DF3E0D01D7E92A5E5AA2E63C822ADCA75681F80CDE87BB3C221A475890FAA6AADD8DC9B45059491A8E2D009AB5ABE14AE3550C3C5962FF5A80B4E89BFB876C00209F5C52318CF82349D6D21AAB1E94ECE569FEB6EB59FF19564A560036BF8B5960D9055A71F8A8E2BC2BC17D00325487ACBAE2F4D29E361B230C2773E68673B239287DF6C2A9EEE2713D6143C7A966E2D22780A924C137B53661F805E77F5517E1A90D541B46238E401AA770D9796BAA8B2DFC197DF0AA81318F27623696D0C5726BE1DC573CBDBD0D019A80C0E48C6CEB8630CBC07C153E9F55B208BAC56E1D3E654B3208313A28357F46C697AAA2C51EBFAC8EDF86167DBBCA3F345E1675BB8AB3CE55F502655FA1CDF13812A103691D828281588AB0F0606FE201CE9A6E818E3C633310F221A31813CBCE44C908F938D77ED5B3A22C2DCE246E01E41B5D8C88EFCC1A2A0F9D59772E8A12FE596E9F47F739163BE4C48CCE02E0D6D14770BF2844B16BD7F028AC367F1B2243EC8CF86D444E5A9764D8172055D6FE7CB23097E4ED60E23C4D88FBF452BE4F18D3CC57CBBDD8DEF8D3772C53B87F36BAB4B644DDA9A64C4D09F20330D8BB4BF5F842C6AA8A80F303D5DDBEB1AB79A6883D557E39F64CFC18EB45B413DF9E8B23D082533A5A0A1FEACD9405648A73A7784C997EE998F0820E524CFC2A2BD050B1A3074F4F31F9D950FB06FD6C3E2534B574ED24E342720B4033125233A4D0FA7D4E7B9D6187812FC99B00B151DF271B9723308A4476AF1D01CDA2554385D9283F90ABCF74EA54291289F1CF430F97A535711F995949EA452B8431D1E0656828DAA3DAADA7F6082F1C8C8CC80A69044E62CD5F0F85A0C7FA0BB8B35F6089A843A03B67685ED89F4D62A2D089E0E8462F6BFC80EE19348254375E8EBC6AFEDDCB0EB4F7AD7E077C454DEF722E60E23A8F6256610DDF2265B183914C15CAB02DF3FB63AC779241DA76C998D9BC7EB72395C866D66541C373142481741B9CED63F9C7F3C8C2D26813E53048A9AD5DA72D8C434FA8EEA0BE8F6BDBCBA74DDFD64DA39E7BB19B88A5024DD6C48FE76D65BFE21DAC0FAB550A87A2345BEBEEBA284C77A0E6549C1AD0C9B3D3D4A47FDD021CEC0A8D60DD506FB70C04D2CF659DE044AF90C5BB989E6CF525088D2A946304466929CB02A19067B8E2FF32A6C20EECFE0E104600D9A8E32880CA3ACBC75D81796FF84DC5D455F0DDBF195AEF3904BE5CF581E0C94D0B8E51B3423F586E77F1A91DCEE74EF33A7D8D8F0EFBC5F7534FF38B18247B2305160923B28B0C7DA8146A6BFDBD6689D83EFA2522B12D6650D3FC0350D38227B7FB677AE2DEAFB8257AFFB5CCD16025A05A63C86431ED5E87D94A6C38A8ADD61C513E565D791BB91780FD64AC7CCD0107FA241AC15452E482A9A16F260B2D79B64950CED1394E51D4F262337E82E7365843195B469E3AB0F641CB3F37D28620396560F5461B677C6BDFBE9D0AF1131C4BC5CCC63E2B0BF3D6FC05D228758D55B2CB16F50F682B23FE4A039541BA7593F35295C5D834CA102CF908EFF9264A35B388C4FC66C1FD1BEB04E0E6CC7799A9DBAF7B74B08099B2D828BD490D94F1E65F16751CFF0C772FC1046AE192A68D928B9850522A335369D73786A1A215AF46D20DEFF2E68015362952A11882C92D64BD3B716076EB9099BEF60D2EBC06800612A5366C2329950F2D3693550CD510F53E6D4DEC45DC43EA7F94EBF85EA8D76E4DDCF121F61C58925941DF475698AF255D9A8B8E7D61DF765A3D98F2B771575C28DA6DC94B8CFFFAC748B8ECCCB28952A0488CF4D6909A13B45A449FBB4F632CF4807D2DF6116CD70F7E28953513EA66680722A3AF70474EAA8D389B837ABF7F12B3DB98811B26C68F13C2A7AC86350870096A61EB57E9B504861C25F7FC1AFB77410AF8EFE37D10851A2D03B36F51ACC1D9D1AB6D644F8E278FA10DE4023A0D44848CD41F1B901BA24DE232122FED32E9F68EA5308B1865DAA7BE19D2534158BC09B64FB80D10AA9490432E877E70D45FA9B74CB4CCDA8045BAF8B33DF6B835EF23415E10A43EFD0FF0AF5BA41D0AE6BBBAC145455C6D0AFCCB1B7AE2F3E69BA7579702D848DD1BA5FE8B8952A11DF6F5150360B21B6C49C36733ACECED593DD17C0C073400E7E451F258BEF69A1429A01EE563303492AB1770066298EC41609DB7A0924CAE40CC940F2DE11624B742CC2EA4ED0834CB3DB527EC0BC47E78ABBC276A80B978B56CAC4BDA9B3D20A991161A108E151A5868E25E8BF73420A078592DFF12DFD7E1A3B746EE35D26026E7918D47DC72E1AAD5C9E01CE1E4B6519618A10E8F948F72C45E2394F60C78BFBEE30368A76FEF69126CC56ACDD2512A764BB10C1C974FA6BEAF043C327D5D2655791575594B8467A863AE456881FAB2EB5E7DA867704AD33E6680F1B8E90134C94F0786FBA8B4A36F57E876272BD7947BE2B688695F8039EA3B7C3A58C60B99BB9C885E5442F875EAC14AF256F8BA2347769E98E99C1CA4002D8FE6470A96FA391DFF45B7A135B6AB2E128E7B0731BDA6F18CD19458EF6B04E9A7C063EE14FF8BF52B14A7B04F47BD7B1A7665FDC20A4467244153940FB89DFFDCA4053FDB74F1E5D9455F5386DB2A73C423086773A9488EC374ACC19EED1950B646957B015436AB70C40FEBE06E98F2379BB8B84A54D182B7214A690D6110C2A56110848D142D42DE3AE716E1815A90C9B02ABFF06BC448736ED24632320B5AEA84222467E182F38B862A53357BD8827E3804FB6A7A757C5C086D966F149E0996CB5ED184CEC2612AB22E6C44960DD60F6FFC9E119BE234EA8000F05A6B8542945A5BBEF3F5E24A3D762C0713C1B5117F750C7D5FEB743DB68CDF0931752230359063E2B6967CCEA18E617A64B28A30E7231E9FE082452A5AA2054E7786EB835DF6C36A015A3229EDB82F2BD5B1630659973AFA6C8972F3BC29673B314ACFA2AB15DDEDAF9B0224B2B1DD8E3F18E552145D3358FF255764BCEED4DC4DD7E786E10857CEBFC2C5DDD045623D686CDFE0BEFE71DC72B981F6F3D78E9599277454FE9A2EA5A0DEB721930927A2E71987811E7EF814CCC3EE4D9B630265341BF86086A392280633F918FF6768BBD43456B6E92B72BADD80B32794CF4703CAC33F6F937B5D0B7EDA498FC3642ACD232CA3B06F4848AFCFE7BEA92442D1CCA44D59CF24C73E9BDFEA20521903F46FE5AC9176C77B9B8E6C8DF758093D2CC3C803D15BFD11E9879A8724215C2CA7EB039247DCB901A28BB29FA80E4CEEAF47288B276BAE83F5ED347D562B937089F7C00654356D4288895AF1D93DCEBA45838314F695621990D33929AC069A8E265D128C131ABCB3D2992935E21E772D1E8A644C08F48C752905D905A5E5CF928C4C551BE9FEF87AB0B2FC3962BB742EC814265640520B4C984F3274CC44BCF424B4AA571AEB1DA456A63949B9DD9259B91ABFF1B484246783CC0BF7F9FEAAB21A0FF4C080E7E07314D0FABAD2852A0A8755F5391D2654B8E95FC946A84A406ED1B0C22F29CFF184BD9078C83408E6657A082629C5EF16F2C7D3C6FC01E2EDFF0D9315AB2B0FA322F35AF7A358668D56A268899FCA3E9F9C6649116E0529ADB5466734BE4B82EC820B2C5FAEA9840E72D59C09F430B42D66F8C922B0DC676936D82CDD73D90FD32F07C6FC4FCF348A8190CCBA0A935654'
		},
		SiggenCaseItem{
			tcid:      7
			deferred:  false
			sk:        '704555B4E5DD1B979A4C3B7A0A0E4EE241D59AE0779CAF0DF58300F21066DDA70C04FABC4FCA7F356AC36C28B99D7A1FCFEF78F38B167CA9D0AB8772910C3945'
			pk:        '0C04FABC4FCA7F356AC36C28B99D7A1FCFEF78F38B167CA9D0AB8772910C3945'
			message:   '0E485811C6F5421891E965C5543BED8CD169FA52C4388CE1A4558F8E130A6F59606D0F027CE6365D922E8C582E65C79C3C75F51E98B9701E4BD5F7FD52D5471E41932B1BD82A02C787930C3456D7B69C52E2635A28B0EC8B89E72D7EADBEF09E62E230E401197FA0D01DCF8545F9057853A5BB4374AA0071782C3557CBD3E55718512E5B500A410E25D805292264B8BF3EF951921508F0913E80EF4227A479D547F1EAFDB94472A537D04B643B3FF2676F5DFB45A82C48024FE79FC3B078DF713C406814CC271D3A3EFABE5E0B3F79DE449FBB0715B616B006B625D67EB0A0F62F57A4B41D36072A6410FBBEDC4FB975BE1E73506F0EC8E1F5864BD352814A39B99BADC5B437FCB7F02B15DD970B36528A7858C9EA5991DC1C59EB1AEEF7557AEE92CA13A143ED16E75EAA01EAE53BE1A139CBA8FB39CC83AE4E09A24DE4159B2C00C3D2ECD88B55205402B6DD3F2B25FB39FF0493827AB265B6EB2D990E6AEA148841160B371AA03D5E2A76EB323A997BA2B0B7CE2A236D16CE090778C9B44BCAEEE818D9A7C8ACF0CD2EB7EF90806FBD63F64E5934D8FDA11ABDD3E30B6E6C1519076CA1F8FC72F009ECA727C587D3A1ED12E635CA65D15A8A11D519B9B6DD75567C7664225CD0492C18BF053387B2F0D78C99E8E3C291906B8EFEC9469F09C8F1DAAF7777AB2E86FBC9F85CF63CE988DA1CB9C27FCE5005F3EE0F51E3CB132574B5421C108C0C904F18B733C8857F7BE0E29459C47D7E34F7C003843B7D9FB2FCC0E175B7C96B6E767D3FFD0347C6F6724BCF837D10E5552AFAE67CFA820E8E15BA7A8E7BF2C6AF65126AAAD2A92EDD3CFE064A0CB56D774F5C677E78D080E02812A6322502F57995DB38EB8735B292795E4C7B6236A1BCEDA090706B5C8A9DFDF1DF853BA73C887A6981AD715A17DFCDD3DA036E7ED20797E2DA618B6FE21789AA459F1580655462BAFA353E389FC7021CDF4E7314474391F405A1FC9E43749EBFE6102119FCAD214E18B5C164FC9D84D600CFE381D670BA67B9112E86A27A70BB993BD6239D02EBC3CF4A8502AA4B0533289E18B43037FABD33BF1CE771F0989DB86CAF02D0AC74198313B9D12DEE26D6F89F773B172827483DA6CF121B6ED7881CB2F1D121FED2A0DA30DD5880376303D138554879B550A93DD100A34C4E49606B390991F2F80E4DE8F1F067D265193D4A1C6165CE43C22644E4C92F4CBB91CA97B0BD9975AE20339D248B3BDB948E06004C5EDE19E11029D37E3F122BAB72732CCCFB606B1A89A9FA7B46DF6C95A484F6F5DBBE2EBE96931128B4FE571AAEE304F7D0801884FCDC0A8D9CB0742151877D972DD98F766BFD4C13E567F69336972BBB01BE1D211B24CF6A359ABCE3A7F690AA928EB2D99F05B6EEA233A9CB46402758941C18E2320F26E0B32E7C21EBEE478F333CD45EF0BFD71AA14F3141058298B1BCA8D1EF86C4E766EDA299761F573DD375AE4EDFF1E400650B9FA61A7513824DA49C7829C1BD3E811BC643F125E2B9476AA65587D03D4D35D193ACC545032C3093BF59D99EA77ACB361E1C3F19D2F9B864EC1EA243160CFE7517D13C88759F38055CC31F9B1D338848999EDD3BC34DA3D0353AE43C328C57DEF4F6D230C364D5FB58036675C9EE9ED05AD4D06EEBF36CEA01FFEC4A9A9009C239E889BC04E21D690DC82E2F37A5CF22857FCC3B4F91C77EB3D713E0CDE2C487329E1B99102350270F20FFB2711FC215E0BA2D5F173B6154829AE0550A2D890C7BA04EFABAAFDDB2DEE476B1E64919932D1D0D57EF3F278199D549EDD62F0C86D1E5FC8AB3EF32EE111D9E3FBCFA2ACB88B68416B35AF2772B02EAEC9EEECF7D2432AB1014A14AB134C1B2E2B7538383C2E7DCA6AC31B97CF6102CFDA166AFC3FF56933F7DECB2655C31476DD7E88857008C534EB2CFD3B77229FCC606A6E37C2E89CB40AA830F15358F7580E92BA6F2D732A485E2DE4DCB963EC28D02E7F4D2B131987DDB608AA411362C009A69F635B6FFAEFB7995ADC707A7A03528214C629010E9DF615DF1862E1D1A8FA655723673EAAE4E4985E29B10FADACDE6B9C22BC6D3560DA06920654DF8815C30BDC2E27487EEEA4C1235E71D8A4981C23F7EAF7A4B4D6838E7BE62D5FB617F6C0026597B9D0D65693C76133C8FF45ECCF661AE78ED5C57163D8082EC5727C325727612E9157723EEF69DD6A263A6B869AABAFDBF87F1E213106FF3C1FC5B06131977E2475E0987F3203669D070678531417E475E3BDC9D55BD71F39C6B4424606D4709E9D8FAE8F218389C2446A085030B5E0620BB735A2260BB4247FBA02BBD5AB070F56A9190479F03D296FFFD10FFB9EF3D96017E11DE3D737B684287F5EBCE9B2256A03EF248F5079FCC519895DB2384CEF18BFA587C0710345CDA854F3ED0242E95D9338488E0C8915AFB18EE71D055ED91C6C60FFC30FB8A24C6D31186619AE540096631101695B79AF788789135FA2FEB0CB1D9B56537FB0B439A1D986388E273AA246C0041F943A07C74342B07CEBEE36B740E440E90657566730A5935330F2BB47F60F4DE9B601AF6E745CAAD617F4EF352CC72B397F30A184B9BA2143988C23EE18D861CB23638E7C2DC019A7DC002151E93BDF64E0D41067CA715D448DDD2E9E0476E63946C8710C2C0C0D9F986BF606FEAF10B71A28650F11B893947FBA883B5FB213D2172FF109F2F98D45D332105E05CCFF06087E502848FD6947D263F5B951E0C1B8CA0BD3FDA519356A40AE0C7AF066086563DA1C217ADDDDEB1DA6232853DDF3DFAD10B41E3252D0149FCB0626E876EDF58C599745C07ED97E1A1650853DD53556D4E4F1EE5B84CEFB1FDC90445BF7F16E2B510D9924C8C49F0F0FA3015DFFF1301F521EE9D5194689E2BC0E851DD88DBD17AE753F1544A8E3DED6F7A21EA1B72E51BE2CE9A5191C909012DDDDAC936606A1C1B3051E52FE4C4BB3F2F1A9D6ACC099BB2883EF3F7ECAB383820390F4A7C1C8A188CB7240D97A421C1923D3C02412167EC244653EA83A8D2555E7DD305854E7C6B1DDF8B33F6BFF8DB28769FBE0197B5F33E9498F987A8F717EB1ACC90804A3832FC3D9AF715A681BC40DB937ABFBE702B0D534FBE8078A9B8D6A0D9777C38B6BCF15F7C71C3C3468E5318723160CEB8C59249C93606299178AE5DBA5C34D4D5B20CF34878830275D68A55E712F1581591FC0E4C52EBC3B03AD70073389AD1E43A2A6489765FB4D3DE9BB4FAB66469792296542D180FFF16956AA82D57E1108B840C4B7B6B7BABE529275B5202581AE2055754492555F086A6CF042244DEFB3AEDB652D0466FD177DF7A820996A6E69A8CED0C521BFE41D7DD92EA3CF28B5FAC30F2F8E8F3A6CF11AA6F47672CCE19910BF7ADA48B2B2CE59F467716807BE727E1AFD7AF37F2913991977E47E4E11D54A86BB8DAB2405C08A22FDA85DF61A829B72B484A22C1FCC4D25FE5E734CE157ACB577729A49E5329F9FA7133B66499777EB215F95BE9AB1F945D79056A5503146391E979D827DCCC25A433CEE190214B65503D37E2780BB5D04F51806B78CE2DC953C4D7AFFEC7BCEAF772679E7C6EE5DEE57E3882CC67276999779FE3C6C4970BD14B5076FF31E389C004499F744E48EE35473010D9FF14A33AD7E0E2507CEE4112DCECC45D1A25168E1282E10B61407A59EF60B506A9E7BE0FAD912547729B42E55501B5C8A1DE95FD37BAC1BD2351CBFC2854EBBED4961391B5663BAF224D49D33F045C2D3CA2AEDB1E899DBD787475E9404794BC6F81EAB12FF16A50B9B387D4783A31993A0C44BC105B40BE48438220B6F563A922C10E719D973A805FBF365E48E601FB942BDEA4F1B67E7DF387496A71C90FF011CFBB7935C6C419B035738ED8334692ADF4EAC5E67479DD3B443762B0EBB6D24D0F928E78AEEF7EF0C5186B93B9C12BEAFA55279C5D00A35D33282544B5DEC9A007489A5F308C021B8622E618D71063697C178FB457D996A9F2BF04B10B0413AB3142A41D2BA801890A7E76F3A9951D38D93149C88AFBE2AB65C50832160C9AFC1590AEF4493D9BC5E01AB03A85FB6EFAF11BBEA601283BE036ED5AC66DE1A4BAB8FCEE18900E5397D74AF1C6DB1999C08B7514BAC753F804A83E029CD57210D1E08B531FBBFA7006D585FAFA2CE41E388A2F397EB384450C1BAA120014281DD2451EAAFA5224F0C4F4C73E0C5F14AFBB3F17C5F24555EF8B85A543ACBF64CD1492590FDC9F5E504F227ED4A20FCBB15F56D164E23CAF2B54FA4A58A2731243C8694ED71173058DA3F902A271AAE9D5DD48B7BE022D3762696B82E12C014A51C4EF7E8BE5A8F91615D491199F1997D7DB775AECC5D73247F534800A8A1B613513A1BB0881C54D37347D9634742C97EA750DFD8E375DF380F7005032E02E93AC09064637030CE4D905914AB9572A48456760391EC76A3C59D8BE15669E52C97F36EE5EBC72FE4AAF2BC5F873B7CC3E0C67EE85A9AECA9A68C3B8354EBC109EFD0501859636AF34EC0AE7E861D2FF110E0CD1763C50CE81BC84956CA6EB55971426CA73C9DB4BDDDD2BD5782F861EFD305E21A35324C5C878CB61E2148D60C182176F80CF2F7030B0259B0118474C1D67A9FA06ADD7AE83A79AA3390BFB02782DEDC07CA485A72A65CE7B02A86C631B056CDE17068DAF43941406775AD5FE2B27436E7C63518A45C101945D1A4298AE12FD0F0A272ABC9C6923CE2ECB682BF92B9645401A751914770541C22919666243D2E085CF2AC16C8389F17C66014A03C4BD7681A5DB80F283DF35E89640255BA03530166BEFB7A217EA1B9B679CF3ACEED8034F75079773E84B7586CDD9579F2459195AAD39DBC70DEC893D4E683DF86502C1EEDF4AB5B98FDE4F47B6C48FA1286A03A59459AFAFC6E3992AC1275137932C4B5C7A7F0928FFADB35DE9A2AAA6174B64A0A0D124B05F3C6DE972B467433B38EA616BA6EC8C0AA477B80A0EEC34CC0CDF296B8C707D8DB602660C14CC7666BE6BD5D777B2F774CF2C114FB16762A379FD3F2BCE01A60EC1D81D9D605C37B5C66A71708FAECA4B0BF76C337E3F65D4A0C7694B813CD02FDC658541FD026B3C608F8E163B026AE249C1689E31827347191B9FCC9997455480AC72FA91130C73969EB6F2867FF03F9402E3C79151DC4E5F17550A7502DB178215962B42FFE52C88F9F00ED1D35E6F2615CE74AFC76916D8B5F97640946D86AD88C5E5EE16556377928EFB68B503598E969FE389889F47FA844197625CBF16F458C3D52CEC05C5F857FD4E0E649B194C5CD3FFAB62DF705EF1D2F4DB4EBB74E19C5F04CE50B661964A4568F9FD39CC791DE51DD1A0B3545C9226E24E9C0F3EC0F64C47311536327AA5A05FB63C0384D42090EB8C7B6B2EE490190583300737A9FBA5FC820DED0A0872993CCF98E47698A91255D3B93965F3CF551E1F3FA413E270F79AB39B2EE77663A5C5E15EFD39AF39452843E9A7A1965897B1F5646EAD387A9BCDD193B0DDD2563F7A5BCFBD8A804A838EEDDC8E7D3DC92E6378003DB6DE00959FE97E8432C73205D167E46AC4BB10B2321A4CAECD19844B55C6770FD727A65FC594799B327D9EDA9BAAA702881FF4DA88D8655D3DC62A1884B001D0A2CDB0796A6D89B996998A98788A74F83209FB579619DD87A111CC4F4E1034BD15166410A3DA0C84768BF46560076E09167929B96D17E607DD535476F100448BFEEA9FE6938A725BC3696E7C20BADBF587BD4F939B33A7B5FCF89B1536D0EEE40715203BFDF5C7660CC4ED15CCE3FF78698B46DFE44CA11F269CDC5BF07E20B17F3A5F20334480CD9D34DF3D53CE52D8548B9457816D1F673654807DC3659AEC0140E41FBB5304FDE2C74D04B4D774A71AA0C08B6A22F2635A1B7438426395EB389314C7756D781417FE7A73D17983AB8CC3E15950D27F1608598C34681BFC5C3A1F7D3782006AFCF9105EEA39FABDE750DD543EC0D00AB6CB97C8DF6A722575E9B36D8E61D488E102A1295A894BAED039F6A78D91E510A8AEDE0C0AE26C9E236BE736E7CBF6DEF76AE524D179B895D7A2AA4C0895905C1F9B39853FCCF2C72673A3131E23507B85FF3D1EEE04ABE2341ED8FDA99211C67E055938477CDD3588D4287C5BECB3B09F54DF195C0E6279D380021C017B9B4EF0FE00D1D4F0CF6519992D517D7F62363BD97944E101C47ED72D2817E1F6CEB525A5FCBD23EE8A1899C01B218D3AA7FB97E413CF31C0F4ECBC23C05E09692534BABA8B247AFA1B4EA9AA05D6ED81A2978C3180072B8970B0CA77B83E3D33C39E9609A22FD2332C17EB3F59A271BF637462FD92CC07BC3D5DEA5D57A712078E024C779550F504951EFD88C369E65B0D221ECA45CB3610162B5A983467512AA0AFA840FD7FE1813FA8C9C9DC1EE797F61FC5A9D2B2B636434AF676D235AC5FE7DAA6AB00DD7AD3CBF07DFC017A5A0CA12CCDE1C73904465AA91D7752AD72BCA4CB43362B89C4C4008CE3D7F810DF60C2492345F1512A2A11D134C5A17A5FAEC8760DE1DA1C56C572BF32F16316178F6EBEF2B15C3B32B1AC1D53814F3783327D47ED10A04D1FB4FB7F812402D748645283FD25ACDDF6B587AD2FF9D05145F3E434C8AC7A6A136BE39F8F52F1B95EDB1723D2942B686746F3687BB3B902538AD272DE61B25F882518288D1423E91E0260E8FC24DB1765C3967B0B038F2B9371B3B23B0FBCBFC41347AEAC912BFDC1FF6B0BDF4D74063C0D819A217773D0D3C4B9B912E4E88A0D4036702B1825E75EB7F27FD362F04D2BC5972499C9FFFA8472C6D1788AB5B37E3F6DD09A9FCCD4311A642071F84399963243C89867C97B10D010F7EC5702C2D8637717FC877F6F8D308B62440FCB956AB2287B4C8E17F6566A571A0E5A04BD7DA9303C8DAE4BBEAD9056B05D20E567EB1F52F014806B09A005C548452DFFE4E0E9832A77B7B4BDA33CFBB797B8FC1CB29D470E3FE5A601D3A8F3426BEFFBA848EE685A3C9704332D92D5BA813EB19447313741D547D24943BFC27CEAE14F79F77CF6494C444DE9DE1D55112EEAC09524DE23BB68F2243E38B49E8A81E35182A304A442D4D6726BEC9F33FA860AFEE24A435F3C64F37D9CBECA20BFAF3A891218DB'
			context:   ''
			hashalg:   'none'
			signature: '8640FE92D4E79AED24513955CDD0D30C527688A9D878F6D0C6E114CA62C473383C162FF7041E10BC90B0240237BCB21836C956D6AE569DF0CD1871BCB19AB0046F8457CA4F826F4DD21CD93D61A824003F94785B0A59F3ABDABC3A316EE77ABF7551A6FDA8404ED9577FD0D22A33221CB86D0C89327514729E9F335B4DEA015B730D0680C8BA84A5B5AAA2F0B839E061E2853DB793CCD5E57CC74CE6448C8AE68CAB16C77710F223379A9AC40EA41CB94C8733C9F13D237F66D2C2A5FF15A5D43ADCD430081C4397961C4F5739E143D76B0C2AA676556638CCF856D25211356C39A6700BB0F70F4567BCAB9C6B001C55569F8B20AC220EC871C05A18960BE76A3E5B8F0834214C11E3B25868132019E7FD34CD0E8BF7B5458229487A04A481A75324F8614CDB160110F6E204B327697A358EECFAEE465B72ED368F6891791D666D207B2EB4625D084126E5A8764137643BF35EB5B61B735E97A5B06CAD2E5D7EFAB9BC6AE66496AE9EB526F755BABFF150E5721E528286B27A3C0DAB74B7A09442A7CE71E71D368BFACC0F27427B38A45B9421CA86BF90A0AE53F5028DF0485FB3654A1214CA0A2A4BF89DF81B7CD3FC0CC15DA65569334F65E217A44E6831AD9003BE9EB8D37A6B250CFD19C638327DB1E28A2C184520735E926D3D615821865D5AE63C75C7ECD5ED6FBA61087F6538FD8FDC6E77FE71D185DDAC08C85649AF258DC4EA4A3FF00BB5DDFE20C6AFDA1F901948D359B1E74DDAC12BC604ED7F3385DB8EDAB2350466B72668657412D5E4A3D76378DCBD6DE4D811BB6342E8082EA26FD7C78A5F74869C66D5861F132F87495690C6267DE456F58D80421CA5D755E00C9F11F3F03D524F7ABC27D5F1A4A156B77B7EDEF90AB2B1706653EEEECAB98CEC87C2ACF71214A0083D7777B4FE7F3DFC283CB574A47C4EF945C053D68181DB0411059D1EC58A0B67BFE3AE05E7144102AEA00DBE3F61E98BF5187DC511D7DB14B0B3FA15CC57F87CD8B82910ADED794679FA3C787E0BDA8FB36B9B75F69A650B55F9648DBC64A918F5CAC3CF818985F1BCC51168964F80BFD31D854CF3A5ED96D03FF2AB666B2B79034DE1153DE52CE835A5D2FAD5EEDAB78F9C5C99D7304EF81C1BA3D3F4855661EAE4AE8D24F72CA44A164A1B25CB362444E7789C0144D0A42D586EC76F402BC47A577661D5A4C841388FDBFE6D1DD8F0635A7F58BDCCAED437846729CA5E89CC715038EE5E553CFFA3D945639E73685BF3A00AD69FF049CA8BDFB1DFD28E1FBD3508137CDF74475AEBBC60830ABAF1869B3DC50A8BD394F118A6160C2DEE09B250FF042FEA3644585EBAA7A259B2014C4049D44DBBA709D9E1417FE38BE073810ADD66CFFE937E43808C497591B5DCA3A0815843B96F2893991B0B614B53B7B5B2CC2B17309DF73F4626E76671B924FB1CDF2466CCE372E9489A9D120B5C50BB35773470EEF2FD4CA05DF9885F1DEAA42D60108C6C48DD32509B6A57DC44F1A37F8163CB3DF963BCA3120237C34DA7709F216F3BD438C256FF909E493F6D9B59D242188319784B15E408EB20F9C606847558C632572A86CE8B8F019E244A417F4F2E801BEC25C5A71E53C5605AB4DC686CD7C37D5FFE55B20A5E3B6C7B4E8436276D4C66DD60CD696E0FCA795123FC1DC27B92FBEDFBB8FD52D6410CC9B3A8DF20B71EC60ED37DAD357B976F6CFD00D5D4D4DDF74E16AC7B25B4F51224B1721FE53F9F103059BA561EC542BCAFA11857FF53734DF626878EB6F966AF5EC3E8EC9B5E963BAA218E48752658B7784AE66E1A77FDD748D344CD5E3C59B986FA3DAC5202BB4C87197F26719A490270238597C43DA775CE059A22C684DD4A64DAF32FBB51644C353B7678D8A81BDBE6CD160A8CC15AEA602BC58C81799A52B48984F6B12ADB84CB7F3025A76F2516F7571B839FB4B514752D3827E36045441C0801BD587859B0BFB389105D25D5521563BA5ABEA48BD515B12B34074223FBEACFE94AB264F96D5B248DBCE17984CAA449AAFE4C69A3809A5A70A486CEE10A40A8C6664A61B51BEAC9C51D4A533C99ACEE542A99297D10116639F453BCAA73D9396E15E521F3CA942E2254D4EE41350A78F2D4ECE26B2B8BFA2ED95508476359C1DCD84D570CA88E42188F37C2402ACB900D8654DDB1AD4EBCC805434249D46FA38609AC5BB15147BC562F2AED6D98924266C14064C07978A435DCD85570E8E6F2ED9284AF63D071CAF77D4BD2A44B8330C8FA859508711D8C814669822BCD6271799BA8C47793BE48343CC8CB9DC13728CEB9A0F0F76A4BB8D0DBD91115BA1C7CBA7FC303347DB5C7802201D6B4A837DEA71505539D69AE1D9F663B1ADAC79A0721800F32D2587A544C61D679E740785F47179688220D7CBED462418CC254E498BC2012D2A68A9041B670CC8BABBEFAC785C63B4639E9D8BA4F74D1FC64BFBE8485786690AC49959431C6E900B9E0680F8C950FDDE96F6E608A440E1B1E14CD997BA7EABFA654E921E3561F10A4A1C0C6BF6238EEA3ECBBD541F49844CF07C1B7A5E6AF1620500F725C76714C3A708F34B51779A45E684BE8E92E2EACF2DEC9D38B6C349AA15C120B9A1490C0DA034F9E6B3094EBC8A6A2467C2D24C0843B21131D671AC6038FAF2EAACB4C1DC3AF8A62D7A7923A52E2FA92AB1C21594A9B3F6EEB4253084726AEF999EBB06EF8E5D053DEEF0E69668E624A249B7F714B822379955CCBC8773C04FE230B0E88FE3598F64DF291E280ECBDF32DD1F61F43876A98400DF1C8FC6DFD43CFD53AA8A9E3E0E9E4F0F1BEAF3E3CA60B53CF528193C15E3A97DD005EC2E16B54C0F1ABDF85FE948EC64944695D12B37D1948AB1A2006F77DBFDB3030AA6FC492A56717F62E5C5A119D779390D4226A5DC9784A8B4821086C7083C99B1DF1CE3C3A98C6C8716D1C55254603D6E6BDE96636EB347EB15871A4987260D3FFA85E9954F074039EEC016C194F442D8258A97E9E875A6623FF512177718812F810B0832BD7C45C7937402FD90F5E5DA8D40D1A0D6CE2ED3707E970194ED1CC8BA92EE86792D498BD9332E58758ED7CFD2524CD3C57A6713A54AD81C7AA008AD675827AEB627717CCC1BF7AA5F7C0B94FF577D39415FBA3918D42CAF781BF40C352AE486AAAA61791EC765B4897B7191EED9916CCEAF7EB59F09DAC54D00238206A44912CACF748D3D2B653F3FDBBE1D7757C5638872F1224BC49C689CD8C1F30A89BB544715FD8B77C01A762FE20AB4254A4DA9101E86C14B76BAEF7D776EF7901B9BFE5F1FD6448E6BCDB772DE1703C6F1D5B7D22D2F9B96074E3680DC5996D8A19F1D2EF6EA4C8CAFEB8D76EC0CEB8075DE001AF35209D3260CE81F739455A9CE933310B3519775275E2C30E94DEC8EBE84828C3D9EC88CE6A6BA76184AD0B2348DBF06C50A9142FD28037D851E7E51F33067DEE3EE7CD8A3FE6738BAABCF21899B1B54A6D88D2118B4DCE566F18F4A61F6F4FA0F201402AAD71B2DD404BED7D403507EB2C917A04F086EB4B71E0DBECF9DE6EAA462EECBECA3CA102E8833FDD6C7D97FBF5792231BDB14A01301A895AFE72175EAE5E50763F4B6C3BF6691247F4866C4DBBE2F77C1661BF5B880DB08968C1CE6D5DD7CDBA7B682EDC5299BE4934DBDD5D27FD9D4760DE5FAC21E3C8E7E45E4C90B068C3F996CCDFF9AD5B2995FF5D80B9B44664DCD1C37C03CC79F28374BE0ACA53FEFB21C59EB76C50A5457707C2A8E9807049C470AA6CAB3AA22188238C24C21D8141481307298B6F559E4992C0F0B9A407716E04D33A95FEAB04AAD4599E70FD23E8FC8759FD28062D8B8A7C427962D92E5413E61E35CFC7BB55E5F451D88DADAD33150B32E65D5A73C9AC6990EFE584D263528450B9BEE689E87C4242326FA744963FBCFC66E1B40763E426BC72C25D4A18DB6A3FB312C9D649476A2A70B3E01DB8DFA501C39E150A0407478F14B18BFEF92626EC7BC2BC8C6CC8FE3A7CFA6312287277569C37C4D03FE6F7F5895E7D6A96DE469BF12D9712882668107F53BB7438F454863916FB8D01662DE3ECF6E88EAEF9EC7A2A1B37B7E2E225FFB98188B2A3328759F830FC65655BB119A086FFFE5EA323DC603C43008603B09E88312AD0867E5DBD3D62A85A2865389CBB40C4C321E4C9363A6A05C0A66351402C5E919D1F16C62BF06B57C38361AD8BD74AFEF92DBB872704F9BD8FEF4D9340F9001FFFE76A332EF6C08703D4877148631FD2EB84EACFCC8A22A73A883133371CC2328FC9C14F7B6B8C396A13A75279BDB33C3D5BD379EFB5C93A990A8219965EE7229C2B587913730F26E153222765FDDB094A4CEFEA11D4C2EFB260736B6EB809C3C35DD1F99B9E9E7593B1FF20AFF832588D5963BA64009E6BFFE7235F12F54763EB7704D6CAB240741B7C7AA51E6FD02D0148E28A9330D432824C57D6AFB1FEAEA0265FF0DD1095E4F418735EED97E3C39853470681F88CCE590407249F84AE1B0F4DB6DFFBB40A9B611099B0970562A32630FF0BB142A6182939F262AF05C94F5D51F4D9BD8003F00C3A5CEBC6F41F2B8C730C6834AE8CC477890A4488A57AD2CD66A6C75FFEFBA93A003D828F490228AB7913674E4B84B9E919ED1045FBA64C7098644F6477E68F9C085B9347C66E27F53FC32B6084AE7C8729643DA8C022266CB1C0B0DEE09639B86D45E000D86F2A1C17E932C141C2B32D2D32B2812E4C7FA0F99B56701C469845B8447EEBC83C04257943C526CD4547093C40B196CDBADF17657AD3E06680F8C02FB6CA17F2305BE232814CC3B63F97A44F963F2EF5A04C38996416C49A9E0BC87854767FB61A2089142CD6B585C735067351380DCF1B76C0E81903D16BB65E0E2C8431B9D916587D398AB6292A52A5A598DCAF4AA697786E926E265957E76526999891AD36F04A194309B733F6FC4C3EE2CAF981F97160DE42C7C8ABC4A4FC6DF86737BEA529A5DEE3D8B910FD56F4FCCD2FEBF646429DF54CAA8C88363D3C74DB6D1B97CB045633FAE5040422A6BC2FED75812BAB179498D4F3CE491BDE0DFBD92A563E89C830C898774F24E802D445FFF7A7325DD941207940027E390DCCBFD6F1BD03DBD9E13ADC14247A168F42E760F198FBF475224CD609B204459964F5E57683B50897278188C75A2A2B7EE739E28F731A56B537271A3391E078F6D08DDA8AF822C5A21189A5DEE04350B722F1B33126ACD3942223D3103526E7C103031C3E279D09352C1CCDADA1771C59912D4419F682D34B5BA1E81964C3F93F3C6DD1848F28973779224F1C48E86FB5C2E31138EA39F621026FB7D0FED6D96B6FF240CF53B33A56409BEA3F950F26933BF8E8B6670CDCFE19AE29EBC1FBBBA18539B2D980C7ADBA798C5271A38E5C6141C75DD0BDAC95BA864C267027DC7F6CCADC7A5C282C4CE15335D5011FFE208CD18843D78CD7D63CDB58F2462D2E8B1B1E7596376A8872D7AC16092F8415E6C033948AC7B39EDBADC5EE4FB8E763AA3ED9BDDB4451E78DFC54F199FDCB485FE2278339A24695BE5080947BC6E7A0E1865B3DBEBE72D22315144DF71BA12039909E2792AE1800E27817BE863A5D467AC185220243D7A6685840A723A144CE20AD340B2DECCCD009941084ACE0762F54B53375D2A5C2EC427659C06507DEBD7B59E402FE50D11FAA96719CCCFBD19F3EDD2A1C948B30397603EF2F8FAA307CF46DC191A5CE8A068DD474CEBE4433CFE77A62E8DF82937CA7F200139B042BEEAD45A113B22EB0FC4151C2E3E4F286602A8CB850AA90B9E2328E6495559A7DAEB873FDDDC5A8B25C3C89576CF6CCF532E069A5630720F345473695C91338ED7502BA6C73D3BC70F24FA1CA10B3919A1C5BEDC0D9998C6645234C77D7FE330943F7521C882FA3705E4B2297CCBD5420488A6F5DFFCF99C5A952C0B15E10BA666F75318D8F767D45865D9778DEC1846B3CD6A7AD3458364BC680E3EAFB1919BFBED8A5660BF2BF7018F8226066748456D0528586B62BF870D78F4CE2A502E49392D41A4A0FB3A93E72C3F7D8A88A63C9DEBA4630D3C8C907B2DB70804C6AB523D99239ADD3472BBE72C98A96B1BB3242B75EA9E4ACA3F178B27E3939DEA24EC5028BC250EE17EC882B22A7BCA45A27A21C14D183170E1EA299BECF1E5E2D2027130C5C18813B95B6DCC22A3C37EA3CA22F2C198F33883EF54D4A44A34C5F946DDFB54061BD854A7F4AE56FBB638E91662A14E6ABE60EF33E08BD5E20F182702653B677EA5E436638B77118B99EF157C22DB8D1715C83F0F1071A939C0396D88352FB90F88FB2C4CEC97E26219F8BC23D5CAE229CC67379961B4AFF2F5867871DCA491A1841C00C011F2D45358D12E34AF38D36ECFC2BDD73E64C3F2367F8558F178AE60A39572CC1890784D45CED174F81E7CB7CDC6B869CD7ADAB95F30B4165D910A573DA37310AFCC683AA4E4C29B102D8D14B7A218D840ECDEB48B947F58EFE02992FBFF83CA50BD1F001390524FE1062317AE2D1C1AEECFF66FB5C06AC12CCC9E0696CEAA9BBA61F6946F36D229DC18AE91DC30BB1F8162CCCD3F30CA0DF93ED20B9B2EEC8272496C22CCDCB71502350C47831D0F143AA9F4DABB678DC0D746CDBC3CB5C3DB809E9DBEB91CEBD42005BA51C3E9EF932F6CA0C0A4964385AFEB1E61206E270915224E7D0A1C02A3C82BE28C09CF9A3E327AE5C7922B2290A15DC51C3DC7EC2F4B8207D5112605167A4F8B8498332098D1E962384AF500F461658BC575C587945AEF82E017D264739BA8DFFEB8DD6C5116DA8314F97B9655FBDC49CA0A9082EE7B1347B44A377AFCDB4B1E7E9E77351F4B3F54A22FC1E181A493837655F6561C116A37BE1BB3E0DE4980DE5741CE7A23690E44264A7FDF277344D5F99D0A2BB2963A1D5A8481F171245BAEDF74BA92B6090A48C7473921E7B845D59A93C984E4A4BF626D027CF3FF9B5E902BD2B1845209569714988C4CBEE14BC26BB8B05314DB83BA9C3A1923CF0A36A823C0AEF7C3C066CF72D827A5EEFBA5B7BE614C72615C8284E7184D6BA37546675D482D0A8D17A14B8B98FD9B9E2398CCAA0A865941C678B4D579F023621B750A44B54178D097BA87F464992E0DB5B04F95D39D2AFECA5F3B8F7BF6518B80517EFFFE8CE771C993EBF3284C4977457341F7A9DACBF3F5C58965AD51DADAC129E77F7B5DDCAFB926C84DE37EBF585F3D643BE862C7EAAD5FAD7A9BE65673747D7C40BE9D875C7E152CFA17BDBF582CEB35CA2DAA235CF130C5CCE0EB8EB3C8CF33ACDCBEBEF27263027747FD078C607A98844A84C1C054739AA2FDF533FA126E10257575F872EE1BBFD52B1EB70D17755F3B44C0061E931D51959395F9253ACFE63DFA8AA8C09981BD8A78114BC5B481AF457CDD37B4A8AFCA2CE5F46471B0BED8227E2A59E71F64C60DECB26D7DD012EA8F84A15901ED6B6CE5C7967F90D12EDD923535DDDFD406D90B7127688C9C735F22A0D67FFA5D0D94C3065C45AA394E14BA83B673DA61B20DCF8DD302CD7E2E8DC34AE7B6A20B9B17EA8E3FF5B2CA544EF4D8D49C86CB0C081429CA099F3C9F52112EC5E49FAF62C1E2B2DEA90BC0668D5C57497C66CC41E5D2690ACDC2F3197C7F250DD193341CEAC388599C2C8C739EBD3F70B619DEE5A9F5928078208E489191FCDBD0AA97A2918CD07FF895646B8F3D83F93EB167CD4A66F1C63BE0E13D6B5F9CEF5D7F38A4B200B50B4690732A03B0D8BF2DC6D8B403BAAE95FE0362BFCF4A3BC1723D43EF4E574A270712B99E7FB7404443BF6BD78286236920B28DBC8FF3B5D6CBFEF06161FF98D327105B36C58D2D416A8E305E1BBF1C9478A2282BE06D62195995E3BC86A16234DD9D8C5A1C879DE681DC40290DF526AD544A1A1D00145309D421A5774739FB8EBA18CE4266C018D57E3314000B19179D2D9A4888BEFF0C8345775B7839AB0A8F6A92C33B658E7A03C04E459518ABA55C02421E5880AB889EC4D126082840CD7E1855D38978699032436FE4535B8E855A12FEB02551F5F8FD5E2F5BCD65BC5052BA5A14AB18FFCFBB3BD164F11C10982508D17AB259C3EC4573B9F93EA27DE3F772F9BCC8BB0C5F64DD8D077DD6FDEE0FDAB0CD16E9BAE5AF9ABBC189FD53AF55C26819542A5CE22ECF3BD769E6DA4EA6E0E160B0CA0AEB942967DE0F92C1598C9B9ED9FAF7210FF715C5085C2DD21AF912E770719BB8B31286A8A03105FC1FB5AF17F5CFF200849B445CBD36423F6C0B6B0366DDCC47B81D94B047A710A44064916162BABE8573D3B713529E736BE3B9E6D4A6C987F4440F58E572EA90BDA23F67E909ACC5D4BDD3FBBC641ABE08BFB47553C9E5E2E501B5B5DAAA0E5524636E65D527419087D49760EC06E61D450E8C562A57BE8B0789D62B678221886D5A116F5389343DA584B4579EBD488AC17741B4BA4D8D731C91D01EA65D9C254437FA4694DEE95EBF5D7963155BB775507026371A4F6BBA27399312CF6EEA17325ACFE392BC58EB6F04B220B0CAF58A5F2E923FBC33F3DE03DD3B9C1EB1D78E9E4D397686D6B77680BC2BF70FB69D8E62A880A00D6880B0C955B805F86491F4BC7C4D3392397A07150857A6D859B9316097155BE5F2044CB1B8EAE97BDC81FE4285BE84160F436C8768EBABF51C4835515CE269D848E2BCAA6963C66B026229AA5CF5854D1FD8CB7B5E5DDE7189B88169DC082F07E25CAAC7AF290E0669FA4A95FE999552AC9B92311B902DD8CC3192B6B7148726A1324FADC49C342F5594DF3E743B98877A0154B34F125A28FAFDB4516E6931359963978BA3F5D9D3255B7DDBDDE6898F8175EA92FC450AE03E527FB12FDB4E1789D37DDA9135E70B3B1E8EAFE44FDC6E6704DCF1C43C048E902B33883E0477066F5D5B1D9F77DE80C94F05E60DEA0D153DD69E38F5AF366D231390446A1400BCFFEDC42B54142ED54B9DC011097FAC01AC0D4A2C76CF4B8D7FD66129E78C188E62D3B15840B4F095A6A7C06D6F033FA9D2654DCAA4873AC74B6C1E3EE2111D9D39095EC5C12A64CD65EAAB9D7B74A018C012FEBE85F5F1B0F734D2B43447E05ED3E1577FE35D8AFE89C70A534E6F2D1A6AC2C41ADE67ED4738D77BE13C0C1AFE9E1C783122AA649E7F1C5A5EC11EF3BBB9F01948C7E9607D0A278438FBEF5245044072E11FC6244C69E84B5FCCDDF5826F6412B07AA489BA4E24D3EBA4A3EDF246A11EC45773F86534BC8E282EFF063F4DEF7D77F7002BB2A24DD1ED5F86465A8F6FA169D06E38C928D2978842F44FE2037E225567881B78131D40096C3BB05C4DA6DFC18134D44BFB5BFF925FFB0820164BDB946C55E9E42293ABABDC77BBDB4F86E324303C5774A22EBE6EFB998D8BA148F2899B589B745DE3DD33FAE37802C92A9D4D7F4FEFA0D79521E9593F90A6195432E43DD434B54109E178D5FEC9E8458FEFB112382521334AAFE212DDFA96B5D1020E658DC6887B64B8201F3CFBB92126C563EBBBBE5BF90AD56A9535F980D40C9D065B4CE28E53E543D2303BB2A87D2BFF24404E6852DBB4B2755653D6EDB1D5FB315ECCD35720A6D61111109DACF47A3C9D68837E14A4F245374D8F72B042668415F110D3C078B8E24B4C8052364535595C7905CD5631DB5CE784316433B010BBC0F7D54D53D1B4542ED6B8A2C6636A31D2C0BC680C287B902BB1B35FF146DE9AAD6429BA24622CC535C45E58EBE34DEEC255EB219A619E21A62C792289189FE6BA80B89797EB3486C679E1B51084AF998849DF9E692EA6CDDB3D64CDB0637A5DF5D4DBF7AB3787621D0E78F19C60BED44B9058BC06F22DAED5B789252C4A6CF63007457622881D20BA3914B162E7C89D55F431B3E95546F34A8964AD07B96306697D6C877DAE29A854761201737D903AB6533FA0F2A9C03146228FE97A32DCFE1C607A0EBAC5A059E7547AAEB84D17191BAAEED7CEEF406F3A95527DCE765DEA77E6081A94B377E74AA5FBDDE4B9F91606CF7AB8D6DB67D5FA14E451848125634AC0B8582EA42FC03CF31E224AAB9D7D1472E000275C0079A11D3E2AE6B39E392CF857AADD04E4DDDEA5DEF646EA96ACAEC83B320D0B273485EE7A20C03051B26EBF1632F5A98C19FFAADBCDE2172477166FFEAE317FEEC5EB853770F7C251CA7B4BD953BFD74765E7A8693982EDB6653C32B85D553918008AB16EF59BCC74C3D7A23FA650D7713B24D31A6117973EF6E0E6EC55E92CE981EB668F7FE3FD577CA3B46CCAD6D94BD272A7F3A64917AB30738C263348C5FE24E8C766138D7D426AD2B390C1171314F7FBA26F1503E43342DDE11D1F83CAE10EEB9A2C609F9D5B3130F7E8D1DA69BA531B6CDF53F53C4FD28BC5698249FC5483C6A15429628FB1F5BB3324EB9F2E1D22F6F5B20FDE4C8CA7E3D2931D5147C17A5DAA0126ECC1CC0EB7D6368DA7E5840919DAEAB048E160B9C19A7BAB56D26CD168974729A98F259BAF2977528FB9A925264418A3542D3D9B188F375A8BBF000620B7C5728148735439F2681C995D9E8E9A0D3116704B3EFA661C176754D828C4BB2D33FB640BD24BCA64FFB7193D2E214F7C1F152CFF4B06BAB728EBD4DDEE5CED2234F66DA7E3F9588C70988D8FEA88FA06219BC49299C561AEFD46C9C81293650EF77637E09210171C00B72FFCA1D56C4CFA71F76A022F42BD43B88B8008FF636C56508492F8C5A7EBAB3F18639614A1ADD31F225B70A7FA48AAE1358A4905F1DB3B6B08E57C09CAE22FEB15501BD62074AE50FB36231CF1911C95D378B0A127A8D7649D90D0B9DBFC6A3859F2FF2F71B3EE5E6ACF32E55B3C3B139AB84D3FD00A213260DB4B1E673F3CB5DCB4C151D60BDDDFAE4BBA312532C5058C36AF46A9833DAC552636166921EFCD0F78F2040EFF91CDE9C0FBDB1EC604D1FD91A411B92FDD9E1DD84491A55A293E72CDC817F19CCBCE453C1F19BB56F81475F7C9931B1EC04AF1764E87AAC3806946251F3CF8DF68E901EBE2ABE271CB57199D2CBF332F489375C949F9DE6660F685C023759132A50A6D0B52D230B71C9091CF7A827BDE1F37BC07C7DBAA6327CDB0053653C7031CBAF92F0822A65345A9ED3CE4F3A5F49C9E58224B20913D0FBF3E6E136FBBE77FFF24C30C2844AC35C15B8CA12CCBE887C3FB7A29331047D1C6F6819E33108D7F46D668DC318DC2375A45F86C6E0BB4D622E9B822ECEBB591B5137A10299311150F08C8964E797F2E9F0A9024A4183F011A39088FDCF95EC97CBD7EF467BAAB483F1946D272E93836F938110362279EDDB18FE8BF30575E73F25C0528E625DA5A990EC01EC500377F933097D9885FA3C698CBDF138566280A35A6EFF27E902AA70D36F9F342A2EF366B4C04CE2F19D42B102057AD5A0EEE936616AF3F62BFA6BAF44F1B73F8824816573FD80AAE346F6F41638DD557AB3CC7540CE3389A146AE380E0960EBFEE6D9842C46184789B11DE9E95E30015C2B2D0D2D546A697D523D1AAD74D8441E7FCFFC0FD52ED017B6E25863CCE034A58532E0D2FFB9993372295A4438A0FB43265F1FC0A8FA4B3C09C663DFFCA8C165F9D7E30BF4EEB545143A0385BB8A7DEC425EAFE8EB129A280390F94BBFE6BBAEF59DAABD8275F5BDE753A28965AC7908DCFF547BCA3CEF96AF385D02484ADE6903E359B1CF531CCA5B4FA6AF13D101E0DEBFB6130FD85E59A1392A62DB04171A6A087A99F7E2B8322944F5F0A454EE487B4C8520D9F29D909411808C702978EC89E16E772B53812276DBF7AC842837F109B09F3E74D1534670EACDBE9DF75CE9DF81034402A987E25A23EABCF3CCFA5BED380CA2B953B31D003C6F6BF4509D926F8A07B1105D748D7371D73EC3CFEBA8032F94B4D0922D70ADF2938FD22F838D5A0899406F012EA566AC4B6B341B00BB32DDF297197A790F376163AE3EBB74A0DDC88D52721F8F4EA76C5BB40548056E1688884B474E427D99E158F5B7441721DF6C734382EBBAC41326D2393F5B2D6B51C71FD1B30AF0DC0B06CE47675DFC30B0A2C6C2132607EBF858D12ED7B38D59C98A6A9963A6FB77CCA77DE8673EB251DBA18C1951F7E419EF632670153E095C60150CE19F479287150187CCC48D823F108CA3EE1ADA2BA5151F2429C33B2E5199DA409AFD011A7C9D9F00B923EB4EACA9DA67840AAC71C0370ED37C2C6DB6789578647687292AE72511AA416357F2B408669C86C3E25D4417F4F520ABA7C97569AAEC3E19B8E73A227D2B50414B6DDF34BA2E3A2D3C209AEA8AEA8E5B11FBC72A940E10C496298B149A3DBF3670028DAECBC30D5FEDFF914187E1EB26B6A9DA4D0B8507ECF62F6D7EFFB325D6FBB6EEE1027672BF0F07CC758CCA75DAC6514CE0F2BC11182BA82E5FD5FE20EE48A7B02AC401856A338C3362FA02F175FB364B563102119FA5BD2F90108F9C4A94308A7A849572898F7A5AFCC91C5D94643E811ECB3A39013CD51C1B7027138BAE0A4ABCC1F9CC4333019E41D3C5CC2C1A76110EBA10CBAF50905EE671E7D2AE9625302ADF884CD19EAED972CBDEB91C9229FBA502B159BFD24161C7F369C95924CB13FA6CF0E6195FD2B1EC4EBB11CA63646831F19C15B36DC4FBB66CE8FFAEC3F4599B2CB41FD441761049D4B6DB623FF154AFE5FAFDAF92A7C5A2A7C0B918B85E47240036E8649F3B7CC375195B06D48B1FE4DDBAB09D9739A988849ED976BA358B0FBD5FAEE462C6E142F1FFE735B27A3F61C7F48F9643DD73E94AE5F5B5BF8A7C491B25A697E4C6174731CFC2242591DC712D4B2FFE6690AB9A516869AB075FD7F5FB3ECBAA3EBBC047ACA7B28C8FE1FCE3C08313C4451B4ADE50195EE2D2A32F7F21434C199781DAA37EC3C7BD26E9B477BE59B23D008FA9CDC0AB4BCC448BE2C148EFE961BD699F59E2CFD512210D67D817364013293E5B50A4FB4B13C466CA50F3308694669452322406C85A63F3CED2885857249199BBD121878B321CB91358D2E996B6ACF47CE73D7DB469BFFA25C96C40B891D56C202A3F32B44BF99E162BCB5F357EE6C4CA7998757631FAB4627C7D1E39496BB92CF7AF520CC5405A3F6793D44BEB988BB172E2DFF5963643EDFA3066F89271E38BBCA45E714D7374B242427E416E507AA2CA12DF24BBF1E0ABF053EE39070563184B6C8CC189059D3F7C08008EF58BCC7852139BD299CFC5161D1D082432FB4371D71FC42D0BA3A99763898E93C3BE5A665A3AB1A214D55A03B7495DCB7A72D0CA29743C2402CE64692BC26DE77B8788CF7C5381B1BAA0FEB6BA9F7DDA14F093722CC528A333F24391CD529AB186E9297EF46CC7237109AC277ED19D20890CF26B92620FDB03F2910D79BD20C2F7A75FDF56EA8AF9BE3B072314750F38571F2CD2293C1FA552677688EC8764F7E655C709EC66F987E6BC85EF60E18FB19297291C2CE94265DD676F9E782ED716E0F5CCF3610728C8C0BFF027E2354ACC8C9E5B0F9337F51C32043C231A3678D068555ED4EE7A61BD8DB7A30252B5FBCCDFB2502FBDF39146865394D9E03C425FF08E31482F3BDD5391E53F0C92F39B79C82CA65E44F424C3B95C290FD99E60B512821ED0216CB714214928D02868CD606238093BD6404F18175B6BCA214AA6F22B6E5690243B9F6A6C2953C1BFA155EB8A7722B6D368B5ABC32566904D102E3191B9598243497EA415D396F4A80CDD9C079C7DDF086A5E51A9BEB86EF8E0993C21159FD7D930F3E8C1ABCAC43CFF7A9F33018CB44180D3337FCDDE8E193DE2E57E9E8BF39B216CD7F69E792BF36EFF7B299A5724206037CA8206F72BBF80504EC0197548AB63D1CFA8905AC1625D3420B8E476A84C886B509FF45160E2853C5F221FD71363C5D51D3E6D1635FCA43B44F852135725DA8301B4EADC9D0C2A8DB9AE48D2D035BE918A14B63A10157A04F062BC970AE18BA87B7DF169B931D4786593228AFE33C3B3044305EB6AB8368B18AF6B566862BB056A0ADAC46DAC4C274C40132F25E7C6B1FF86C193C943188422D962D2733455D59CA30F62C78C434E0C087BBDF15E1FB3F480C9F9262B89DBCF8147A69C00C20BB2C830A5516795744B2D1BAE141D0FE2774CD4D949C65158A8019C3EA060A6A3A384CE40FEB5ACDB3A047F6CDF99DF3A289AB226AA964101488839598B7A01F81741F28DA81565616F0CD557D696DAC69B8191B12D3DD8BF433906ACF5B5FC6F73B419B6C0EA275F5581F19514BEFC1BEE23897699F9327CEF3AACFAC0B10DC95E6BF1E7A6DE999CAE346AD98F94DBD0335CAE12BFB689266EB7E1D51AEA724DF1B0BDCA68812E97295E67030ACFCE44C8097F6E917BEE8A3954544A547A03D8967102324B85EC98570A3E6CC743FD2E3CCD0A220197B17A9CC079844DCB608D56EACEE18F3C737FEB8FFA0DD99175A60109C9E3B9A46276A59B37E283116960404A033781535AAE733008715EDC5D8ED1914401F59BC3B7B25B41255BC377B131DDBEA25F4C52ADAD0D3BF7531475BD14FA7A1461F5AFF645391E15481CBAE311F0A7B8C12790097E2061B2B7DCD293DFC1BC8D25AE2C958824ACBE3D704A1117AFF9A2EF26871B5A6F07A3A01D587AD4B3E188DD54052EF9D188E529E805BFE1AF731FD6BE79E8B8FF0EB20B34818DCFA1D7DCD5AB0CB858349A05EED81EA1DFF4603C4B1191E4D0C726C42A28A0BC87C18260EBE58E9D2A76337B20B1F5CAA04D532410698E1C2992BB636C78BB8F6868920A251BC125C45E12B636FDB273CA4D4A967700B6519CB770679F9B4BFCB313E45E6B953F190B13757728440E9B4F44197A0EE52D6DE9DD22D0B6499381624DD90455E5A1BF666EAB1D1DD535308C044A55EC5CF5559CBDF7C0B5A9216641FCA6A88A41CC5A27B2FF6910BF96B7D9CE557FA3D6E0340999A03248A5B89970B8ED64799C944B9CB550FB5FA281588F55B04135830A977477416FD0B8ECBEB3F1FE97CBDAA968AF5A6890091D0D2E863406DE200454BC2E65686973D4E8235C8D5627F9DD52F77A72E348D925CFA87B99147ED63DA9F3ECE32685924A8AFF6727403C91EA7642E12D25EBC1989DF905C5C1A4913782A6C371B3C44399F0C3D9459EB0101344C3AFE0C273CEE2A72D1661615CC05DE82B08E8DCDB0EC158D4A490D7A874D3E903270739557DFDB50DC5BA4FAF25460EC5948A300FDCD7D5E12F55619DFBB2F4E7F2628D518F15019771207DFEC95A69FA66934D619A09E1E2FA693E924250C7F084C08F6F1559E8AF9B1E4626BF5167216DF39508F61B906E80919D9ECFE142B2EBF12222E833E23ACB6A9EC10EBA304A800F5D2E3407A021F36644EA0F6D99CB59CA6B03037E0BAF80EA1CEB4621FD1C62AA4972CC0C9CA9C34EF1435062303D6F9B73BA6DECB5FB01ABE01FC6930868BD1B78DF7C97E713C418B67A72260EF1E37401E3546C5D8F317740BAEC4FCFA807534EEA8B40FC24CA26E568B47309F3D1EBC4BB8928B3487B56E08FBBD0415F2CD338D1A8ED1805112C544DB3DBB5CDAA92ACBC0A48683EFBB6EABBE391FD569EA69D96C6458C4B4B7F78770945A3B4E0D554A057BB7BACE329B7D6D32C0F59FEE9855F33C42317C52229325310BAEB68BEE880C04DA44F23DF531FF3F1353DF6BB83F33C63C342CC2C1AD7361300F1BBFD1762A5D670F71E0042DA535A71F28E28A565A93C4CF9EB9A770C3775414F2998B3F70A2A55BB28E0A00B9AF48280F3143BAB7EAC368F135FB2E3922C2ED550C68CB4B21CB00F2410887F24028DDD0B3F2EDADE07C696C09ED51AFDD5363E6F41CC38BD26B9F7265CEA6A868A7D40368812647D69BBEC5366BAFF9C41061C38359E06C102758DAFFADABD750AD1EA7660F8757A0AC943B51B82968C0058139F554149B88AF763EA84BABCC07375DDAA0869BC0CE4A0B7E6D747830B6573CC76BC47C55756223066CC79286BFB1FB968DF3DD64DAAC615C90E06F7589FFEE6B7F65916ACF932C8CFA38F593913BBD25073E4481E85D3A725C10F8D14F8894D5F093103C59CD5444DBDE3456A34172961E186D8869E2B14B0C5D02281B5E19E8B791E5FA94B4A46898A3256322680A233D49F535FE8BD7C22E3D54D07BC0C60A4F4E00AC7D3098F1FC6C28C3F38381CA08A123BA69C56C88BEA8741B2328339582C5B7BFC5DD0F5BE91A2BD4A617F9A2902C9EA189C81B7F30FACB853F4F0F4B8B5FD5FA8678429894BB7FFE4B9AB72F5D42AB54A55A851B50DEB2E59E0E22BF5768D5304A9D14AD71F1DD586AB77F7B369C951270EF7FE4E2EFD63D90E8B4FBE75072CD59EEE1D3DEB38421C7B5AA51EF8340B0890F6DFA36EABCA4DAB67F899B8CF1048BFCA1898EBEAEAB0889BBCDDCD755C7603DF92B9B2362175D05C1A754F9B898F221EF77B4A050A82406C37094F08B72112BBBA414796B9EBFF8EBAC132218D0E5E9D0893F055BDC2BEFB78538CCD4B54243DBA8990DB958138F4771832F48D72FDABED59567D43D5BFC83A70BF3D7F81C4A9ADAF9470E293B03CCFA921990D8CC9E5C06C941C0D2E59B5CD83EFE94ADE51574687ACA5361D2EAAA0D5C04C8CE37BCF254EB1B26B367874F62ED0DA5C44255BFA6E865B7E22F15DD310C2FCF3B64164C7A3CD657C7732A349106D6D95EA56041EA3B692CD3CCFCB5C7A8D7F7104A1E7004881BC934CDB1CA6198B9ECC0793A2D0E9145B06F13E86665CB665E3D1B20113CBCF64D3885C9C950D878135815B5A532DEF703EFB89B86463BC61CA3D0194C4B702E090DE447020A68D04455C009161B362CFC242DEB6D10FACCE51EC124995BE6592FAA229F5D3CD169E26557C43B42F0D9EB6336954634CDAE106869A71202477B5FF6EEB1D40D26A21E221CF14D436BA6F1B0373B390ED0213CAD867C47370FCAFA95630265DBDF12815CCD0782D8CB3933C8B3CCEDC6E88B89E1BAA5606F9D1D844DE90004335D6EC69679CE33EF3D45D6EB9392C19BE204EE4F83015B5EC5426B9B7805641DCE23E67CC9F5CF93183E27BA722AF340111A8656FCE18F6BAEF2C145DF1B58EC111884ED0C66AF949319E6192B085B976350B686812468E929E8CD8E9346B99913C803C19D1005384272AE73E7B53C74B60BBFE6A88603E4CFF9B4A17576D3D3CFF74CEC296F48658B446C0CCB0FB90A33379C9E36A17D9997F4B96FB6C8BAB01DF2D4D2A5B837FA7503B3694F4A06267F5E94A0A4885A98666BDCC75E03F8AA1926203DF1190C4E3A58536902FCC8978E7FF6B16D59F67F87E5C9004C88C52D24F0D2E5906D9522ED73652D289A44A0A4F195D48955E815E044A83892CF2FD3E97F0C82E86931EBF92A1C6B71F115B271C4F08CC939362612274A71350FC013AF6F5987CFDBEDC9A04E02FD0ABC9A2E6FD4C98C008309DAA60E26A9326D52DAA4CD3A496820D9ADE830A4FEF991D1DEA1CCBEA5E35931761E6B47C47F07E051A14A0FD6EA92750466A1CACC8B28208528D7EBCCE6B12289199EB731D6F195D1021860F664FFF5BE8A6F06C78D825CD06077A6A0BC6B25516FCCA46013455C3C02BADFA962B4EB7DFBDC06FE83C22BC08448A494441ED1EA70C9D7D02A5DFCABAFB7C18265E36CA2B779A628075199C37B743B84B9C8612A29C3BA825E2CA20240F6355F932BEE548D380F39BC8403318BC5497F59DA3C4A01EF960BD1F9F8B68445E15449007C0C2DAB59BA33C56FD947F7103EFD345FD65917711AD5C4CB4F85A51689C7A19D85B89ECB65BEA4312792518CAD9BCC88BAAC9228C8A5C869E1C292FA423D8A8CEBA9576B8D86F1811F2599798A61C97F3DC92635A3228F1E27177722E78C69B66F36FD0B92FC76D3EAE653A71F3D07B146A6BD8DBAE275BC0C1580DCF99DDB8F5C01F1C8C1835F8FBBD21CE4DD700E1995DCAEA36E40C2066ED28B70147B84E7F522B87FC6D4DD5DC55803537739DC8ACAE49B6BC345219D220549A72481E7A53A953AA18D09A7044347B8AA8DBACB8E00B4AC140D300FECB4E03C687D0712FE6D18BB901E9B8454DCC358FA7A5A03B8DF924C7B7479EFD344FB91BA5AEB2F434BFAF20B3457D99CF2CE056966B23467EFE5957C866F59B4231F9435F960F6606EA33BB2D91ADBA8EDC4895526F0393DBA08115234E70099E4D4F6D391665797273F6A0A596232D456460D56569B370DB8BFD064072F2E6EFC13D489E5A26862836081EF820E920346BF3D6AA03949C00851BCC142862F47979F90ADD5027CF4E8811C35C9807A9EB276B5E27A7A412D4D1510281BCDE599815AFBF30DD68A26420F7C84A0855450BDE2F52B854BC9307EFC7AF066B03B6C354179279E871F9AB86656409EB0A21AF6DF82549E68E726F3BA624945CA3F566758A8628951423FC1A180E919065C3B03D661460A1FD0D39705AAE0273F820CFC91A419E11F294A7B0DDAD0D33A189E639376E3548F470B0155735D4E6D3B1B7C0F59CCB87B90AE6D4F0F6CE1FCDF90F6D90E387915863BA5E0ABBB90BAF109ECD79E3FB594BA02DCA76E18B54541E1C7541B80AD39991664A999F23C844414F3BFD7027F59AB82E2FB1A591BD1AA645228796585CF93BA822091938B08F62820416DD277B385C50A218DF1836E88E7A5AA1D9837EBB532F14441B94531D143CB1160C76F60AF02FA9FC716D7D9300ADDA1127D26B49EF9E454F18BF427A07C1283A8EC769FE8DB744BC8346ED3C3883BE254DC45499B4BA3CDB2121A8BA3844BC70098DFFADC8931C7F958510B304F196986A88BD6E656D50813085564D2AA47532BAC747C18FBE43F3969EF67B236822906E0EE14D40031F331CC03587873C6712B8F8E9A25F62AE8B0E726335474AC0112422015F496E8A800AB5FE385637A91456077C3CDFD015FEB255054D62B615706F4D3F11AAB55C67F74CB245850DB54D9050789FF3A4DE8DFEBA52CB610D0E0103F63785A5A753161B80D042BCC0C1856BD05777E8180E53BF6D0CD26681ACEC83227433875063F11F2A9ED63A788979EBF3252F1D32D5D6FF348845AD6466650D5FE3600FC8F1FED8D6641DEC3A5456E809A84D597EECD13B05E7A46994C7E4030DACE88166ED595E290AFCA4ED37DE0CFFAE24B9BE6AEBF846A25B23A9F7C3F6DC8A4413B6B586F459ECB8FF711FF8B182EBF797824FBFD58172F39D2CF20ED3296598CE6DF6B874214D625184127480A4ADE2376A05FA6A1DCFB29F948A6665E42EF376284D9BF2F7B91CE8A70B49E5FCFA1D4287285C30ABE4907942DFBCB0FA80BEE784F0DCA0B55C0BC4BD0FC7EB877D64223BA393C6082B36B6C16A626F3B89C4349B6678089D2F9EBBEAB09BD4C46BFFB4F6CDF9D769298B57699384A633714E1757739AB810A0744F7F93CD4BB6D171DEC2FAFEFFD658887C185413C7EE8B0921BECE836572049FAAEF868F285297D4CD08805BA95BCAB87149C62D69C7FFF3BA1BAAF20F4A9BF895ED46BBAF1DD4B097C597DAA224850C9AF75B9560509DE312E84F8A84AF376E7149B1CEED0A2803084BD7E4076F7630328AB2829ED808296AE954DF1898E69F2735C08ED158BF4F5B0C5789F517B40637286FBA62A25D6217A9C7B95EDF8B74ADF0403D21569EA894DC2B01E9E9A4E6AC8D4B68A3D65F70A75C1F5AADB75D04EDDA51DA045F9047BE4F3EA29F86B3B81DE9E859A650F85ED5BE62DFB973B4431790C3228C9D8F600A41B7250BF2E3984C6B706E316928E99BECB3192AA182C4A7C3ABB8FEEDFE3A6101C9604B742482BF0ADCC8FC136D8802401A2EB981E6FB5BF1FD8FA169FDDD63CC21C3B571636C69BD142C5EE3E4B5BCAA88B6C2B73A3474A91715227925E9A7BC649BD94CDC757968DC9C607BB91486946617E3EDE0E463883CD965819D1DB5F38D444CD8A5F7B5F5F3AFC81A3806CEB6629FBCA9549F74E22193A3E856EE4D1C9090145699A8DE2599876DE996F7A42AA56DE11CE830CE888E33A115F6C7CD4FA2CE5AA31AD09749A2EF8B0A8F1F5BDF3E82938CEB236A19DE2CA3647D7995B003FA20BB6D9634075973BA8B6DDD4A5FFB13C792E6EB8843611AC544B8E011296EB9E5FB1004B68993254FDFA6F92F81A7EC7710938F445686F7088FB41B3AEAFA865086EEA4034518103F512EB3790B229AE33ED9B3C1AD706C8DAAC2107EDC487DEF9F08036CF9E6A04555AADC7F8A493E01E923E58C60176288D0198622447E20A8E14E6332937FD03ADDC940842AF577A62371EAF62D5BDFCF7EC37296D9665161F9567A74D46D05CB50580E052E37ECC1C474BD716E9D7D64F43B5DC6C5C2B64D30A8A8142F86B50A0B228BD55A880CB86A60B5D3A45B1DDF50D51ACE968DDFC926B0DE7F33C6724534008D06F980F5C68B08A63A7681164D2A6334BDB0CE4B2433AD747831A3B35C7961A813E61DEBC3588B404A17E4DDF8E3F3E67D1B01EC7FDDFE5B319E8A8CA05BACD0B6A843A912F1CA95F9B4717646C50865BDDB668C743B412F3688C52E8E3CBB92E683E768B9042DFDE2E4B45A39313B6F078424CF030A785FD6C6B170F17D0BED1DB95D99B89BB914EF137ECF025059B2963DC0C5CF3CB55BBE32EC3312950FD660C1F0FC621F7D93B712032A67C293F45D1C28E7DB43D74A0FF64F62B127A0DFCB4CCCBF75F8B298E5AE5DECA101AB7487E52A04EFACF8F2263A8BBFAD20F50739A5A1C3A0CFE7C053E1A4B2DE26235198C968E74A151BEA66DAE65A4339943067700F23B28C4A5E01FCA39B936632832315C5C2A4368E31B8DC72BF86B00D57826271B1E59EA823DC611516AA8C6E722C9508CA00D84B09E55CA55E92692964AF5E91D1400C6295E69ACE1870C4A0C6CF7C52E5886AB7089A5C765B7B7AABB26E71E1DEE32933C1830B4464E4803519152FCEC993CB7A7C122A1E0A8DE7CF3470DCFEF04F7A34327184B2E71A184AB099CB2F67109C346191AAA0074DBF918C58AEAD1028229A236F793E417DAC163631785B5D0CFEEB96BB7B1B3711DC25CB050F8D8B2CA1E54C9EE051BDB24864468370884CE3F9613543F609F6ECE611C98B1C4129D5F74E887717A830291B027B7425FF92D66D6CAD309B94F610B1DAE6F6F737AB303641A8EB397B9B65CF9306637A7F9FFF7419740698EC4B846CA673DDB2E89E694679870D8ACAADE2C422F558047785ADBB20B8FA76097BA9B0DCB6EAC3CE229AEFF90A4B35EA676F3CE96B7A9FDAE4A7830E26803412759EE2919E6467F85CB5DA82D27DC9379041E168119CEAD4551A92106D745E0BA38CE5B9885463FFE880EB6866907BF67DEF9C9CE4F7F1033924FE54D1A39525829C53BFDC14CE712A0797D781CE0E94D7D0B93CB4210EA989418BD464D4D0DC3FAE3A27C9A8FABA770A886D1C7FE29A2FAB43091536742BCD595E6C57C3504F73558C8F53E849053DA6D5130EEA3FBD7FF8F265E7A46A0CA85684530499BADA186880F3382D6E284CBF1B5F540055D093598335D46043F66E5891420FED16982F4C4C1897067564923635F2A64BF61C54F8B6267626FE7575BDB479A5AB0A943AF2757531405D8C242D75EF487DA9C6558E3EC12B0E59B2301C7C3982C967170397A4325BB3F5AF620BCAE624A56F49762542AB28436C8A6CDB8882EE22C4C3B064F4F0259C770649660E72AC6DB3892A29C54CDB5E664404DD3F38DF80AA532D23154E0416BE9FFE15098F86744734597C673B256BF337F8C48C659ED18062717E13916E951FE60B909148A1339803A089E9D061365064E68C6C135D235D3D0AD987E981BB835673D9A51FFD23F26D1A24C1202AF2F4A69AB3A19934C2A6D90E631FB1524236437299D45F68A3A47ADF4CD5393A032935641B619CFB9F48AEB2741680ACD79F7981432DFDDDB99E1EDF9E1F4C1BBB91D158C0BBC4840E0A97D56DE41A7035A9771C38FE62FC7B1E8EB8F1C1CE230D14B4BDD284B18EDA47366180BFF9D41FCEF815FCDE19CEF373A3D50563CD087741CEE9CC59DB2AC8F3810796C792135E94C07A3AA1A7F1EC8F74907FE1768CA82D196C2D07BDE44DABE4A5094D00E7C76A7E2E8BBBC84C8372D12CE7C2B8B1287D76C18BD71B872347152B7D217D06EC8282DCE59592D13A97751D0708B3F78205EBA919278C2C17BFCF92DB33231E49D4439D60D4E3A9C9A7733848D8253041CBFE024BA8578FDF71D6450D7BBDAB8B63F2370F272D20B74EA2F08363FCF1A015F1F55132E8159DD2941585F5292346933A3B82CD27E5C32AAC46416145AF03E4400AF72F84E9B25E5A8D0B6C62B4831DA48F14795F8B57D7D6288220B765EF459CFAF87AB658AF9B9EB502CEC64B0BAEE87E8790E8069FA1979A6B413763217B8E7FC3F52AD32635D4393B2079E707F6259A76BFC58E6F09C8BF172E8125D3E7C338A0D4E53C91570F94FC97E05523518A281BA4893F4FE9CCB13A91568004D8E21853943BF4F2601EE9592B3D2997DB3348F7E01BB47E220B7D2C35841206020892E3E0C0514CA1CBA9BF29FCD0A52EDB2D0535CB1E249236AE116CF178FE7D91A2FCC03861E8FCAADE85018CB4A6380DFEAED2499E45C7381F176C5352623133BF40E03A77F3171C4D76F160CDB87CED9773DEC40B659B038929BB5C19A83B22F349C3FC2C92D53AA1A3B8C85CE40275D7F5FC57B685517E989C8AA545ED146A425BD55705A6253BFFF051D3A37D664D6A4D1C3BBB7FE89589088591960168DED82F6C8F95A7744A1AC2E3557F051597E981989308397C302EA52481710C3C470E05B6608FA6CFF81636418F4D6B297B1273BF2D05912C3B4441A04389E18338A0B2AC8866279C26EF456FD0B2B703EB08EBF2C3E733EA426031747591CCB15B7DFEF67281AFA9EBC97C9675C37C0D5619D94A46862083954AFD948680572E4B830FB3F2D6FC34FCF001944222B5DEF253D8227F11EAD928D9CCCA70296B170D4F59677A2DEEBFC3479DC04E44EE1EF2E33B8A9EBF755B76A744D584C5ABE64D62C70B68C1C5EA283D5784B3344C2C40ECE704F7EF05F355DF20508A506659AA6DC007611C72C7A784AA7ADC93BFD874E57AD80E2FF4E8C8DE8710447CA17010670C5D75EC673695F5CB2C14B7FE12C83CD9AD85CA0D8158FD6ACDE123B2815FBA194EC770491857B16DE9D21F8FAA7FE33F8A2313FCF8ECF893EBF1C90AF6E28239DEBBD340E772FBD4E80BE76D6374E79D8FEF72EF5D8B9ADEF04A7843D2D5B54776C460272A7F4D454AE93323B5D49D428A7CBA9D1F5C2C2D5292CF05A81347E0D7B84D80F014F65F8C186A04480B524104690526D48E562274AA32B106A799E47DB28A745E58F2AE10DDAF3A384A8B62A7CCD436C26D182242F8903A3FB5146D86CFBF8C70BFA7E1C9678A985930B6CF467F71D792A3961C76F2E335D73D86D3C517583635E7BDCA89F0467892BC02ADFE9E4F9ACE506AEF342ABE60E674526652C04939E18A282D97E6E20F5BDDAC6683348205BF9C1C157966419E0795864E398F2794C8BE0ED656AEC28EBB1C0EC724EA12066C95BC34B3BC815451153EB72EB5CD5038BFF23240C5D04465B0D7BB3DBFD5532EBF1E980BE0D61B4714BF0A4E3ED0381CF1858A99D70F85DD458572AA5A63A03BCE530F937BEA00A1274CB7BD333F39590646693C99EA1FE0409E77FAB130728BC060A50843EC2FB03BE69A3095FF517C458B544DF33A103FA23ACA992F039BA5B6969EBA940567FAE110A66BFD16A9246486211A05F5EBBADCE644ADE368E337755A953A455FBDE17C67A37DA6B3D911BF044B9E7A68D842ABEC1F49203ECA854AC5C9BD2F04BC859C1A2F6A41A72BCCFABCFB21474EEECE896057DFE60C0CC48F92CC0FD910A5D07324BC7F8BD9A732F4495031B3F0271ED1AF873D86260EE227852299D76563272A5CD5C91658AF2A5E395090550BAE4392BF48325D362F6CE39E93DF78C2C7E3E58104D02DC4C7165226E5043460C41463A607C627565AF9979EF3C3BE8E81D6611E22C5E340BFC75C68216FCB41A58914AAF537829790AFEFEBFBA5C1A229B47BC4F8D1BA83BFF46BC74D6014B1C5F5FAACBBDD37E2FDC20BAEF1C5C12B0E3E8AB16C7070D2D5271D4D0B6802B6ADBE3D5F17819C7A23D608FF03047AEDC60DD8C29B9C7398B82A9358856BAC6EF70999A822DD84A7DF48B783C52CBEAE6DC69E64607296DAD5AF926323FB659C04C29CAE3B329F1D7572294F5A28BB3D754841881628E0DFE3DB695C3FC75461BD03E1E7F041589272E23B80E445E1F4F43A7143E7C578057B39259D28CB5C718246E63AE35D567DB73F2ACC01986017E35BE5494D4770AD98E143AA'
		},
	]
}
