module pslhdsa

import encoding.hex

struct SigGenTest {
	tcid      int
	kind      string
	iface     string
	sk        string
	addrnd    string
	message   string
	context   string
	hashalg   string
	signature string
}

fn test_slh_sign_internal() ! {
	for item in siggen_samples {
		kind := kind_from_longname(item.kind)!
		c := new_context(kind)
		assert c.id.long_name() == item.kind

		m := hex.decode(item.message)!
		signature := hex.decode(item.signature)!
		addrnd := hex.decode(item.addrnd)!
		sk_bytes := hex.decode(item.sk)!
		assert sk_bytes.len == 4 * c.n

		sk := Sk{
			seed: sk_bytes[0..c.n]
			prf:  sk_bytes[c.n..2 * c.n]

			pk: Pk{
				seed: sk_bytes[2 * c.n..3 * c.n]
				root: sk_bytes[3 * c.n..4 * c.n]
			}
		}
		// slh_sign_internal(c Context, m []u8, sk Sk, addrnd []u8
		sig := slh_sign_internal(c, m, sk, addrnd)!
		dump(sig.len == signature.len)
		dump(sig == signature)
	}
}

const siggen_samples = [
	/*
	SigGenTest{
		tcid:      58
		kind:      'SLH-DSA-SHAKE-128f'
		iface:     'external'
		sk:        'E02DFB4E16F959336B9DE70F9A8BA5FA62958AA179327D8B79C8278A3E7A3ABC9E84F23F025B879A95C868FEE91B41125921D1F337CF1DFC574CDB12FC49DAEB'
		addrnd:    ''
		message:   '8C8361FF301D03326BD745F478AED0449438092A6090F61F3945DC8F854FA0DE9F4BEAD2AF4C08D1769E08ED8DC223F36705D04ADDD57F7755104B39EF79D174C4D2B79BA1384A6482E700DF084C30847ECB0856C365B156E68C0AF9B18BB9767D1139BD47A1BE705C93AF8E2C6504600AFCC4A8F04E85FE90FE3D60A9A6F832762C450CAC3B814374F9A54864425524EDB3A0A9BE2FA3C21DE6F9C9E5336A02DC13D08289F214ABA683D79311A3E48AC8239413A9D44646AECEFEC1E628C64B8DB7EB48CC1D4781C74A7D047652911CA7DFF1AC7FF7BAC75C9C9FD073DBF524884DE6A3BF8C69B9CF130A639CA2E34E9F729CDB4C4E99735BABD535D71695D1AE1AA759A0318F44BB3DFB186A157331D277E708ADA33E2FA787D54FD024F7CB2C757910D4B5C6877B4A7F8B7E40FA30FBA55ACFE1C147272A7B0F67B90A8E3BC87A5965466ED72C46C9CAF4CB69ABB6EE8E595E5FC04586DABF7EABE20C50453E4BF42AF7E8BF5404BA8F264722E7A927F2730950CD86BDA4514E05C3DBE7D6F01116B212D2A86297AA2CE67EE9D729C54286C9E3405755FD07FDA04A57FF30A00D101F4BACECAEBC5749A72384C4A1F2995CC20C87E40030625EFF8165B9E1514F6A428ACAC221059351C74087B85C067E05043950800B509BE90ECEF1410E1E8A2FDBE1CB1FF89D95128C93359B1A712DF0C373D76C802B4B0EAAC260B7181FE4FDDCA2298AF74179DBA5D0AB565F45AC6E850961F21B67D1056BC26171793BE337E994E1C6DFB2FA2466F3D45130B6D00B34D9F3FB57CE91BD69083CF165DFCF7922DB0D3051E0477805B9C1AD253A0DA7B3C65048B50513F7C432A7272B00DD28A1F98C3E5E84D28422A8016AC656F0103068F143077073AF196CB423656A2107248803154B3E10A50A58B928B52C6379550C914C0701B0A50ED77C6E2ADDDDDCD1B6972ACF451CC2B5F845B716818795DBDF004246F2BEBBB2D35A6700C59E5010CFAA3CC23F58564ED83FC5BD6378693F7C34C82DEDAC7BF35A69289C6B9AF5BE031B8EEBC6120FA72E2FF26EB1161CFCF6D39ABA5C532B5E9503D54F00847ECAAE77D37F74601317EF2581180A11F62FB82820E965A335D79A034BDA2AFFCDAF48FD80A745D42417BDFF5E922BC662E1DD004ECD33C6C82F1E19549977D0174EB8ACDE6DF2D33007F554B02DD254F1EF9DC3AA424D855B266B737B76DB1A6B6D2D31E61CB500A488429C528FED33A29A8F30B3E33D447F9EC8936D975B72A347E39D6075EE801F51A6E887CD2324BAD90BD7E97F624E0A8DA7D59DD4514B70CA6976B3A70CAD7178AF153248D227746567BFE2CC3D0DBE97446D235FF9CE67D8305AF5978A2298EDA3268C20E54FFBCA3497A2B824A1245E0E3DC9A49B149F3B361897CDF1A9FC0A77066D616BCCD40E11BE7498099DF0C828E741872C0FF41087F8ECBA5E0C89A930AC5514694C454FC4F6B49024263323D2F6DA7B522DB6CD1BD6ADB11B9905C54F99BF3DC0C3BE026293B4E3DC10E735AA085463D2D842EFE916D8284FA8E278DA91A00C5CDD2C2759AD54941CA0E3F4FFFC5AFE12DF56F0A51B1AECEB17B0B628D083C005E6320406674229C8E80B0303C440FF5F0A495E51A6F28EE1338E9CD71D7C28A4E7B93FFBB9085C3DA89698AAFC1F7AB487D4A4F927A8BE252EBE0FC380D25F80B600233EF48633AF4386FA6418BDA042521CA97CFDDEA40BF73482EDB89FC3A3FAB1689C62CCD13050A2D8CCB3B559B0ABC863447559311E9D860AC5B683511B52AE1A726D4B0BB5601FD62FFD419102F938700ABA16511524D6E86E82315026D1D50E45B853E91CD21E5AC76F55F485F48DF706A923F160F3D2C65767DDD4BBE64585F2C6868FF13F1A2DAC7644E8EA2D504B56ED366B56C7D5CB48442937FFCAD10B574021D540E4E43D157AB835BE1B0B809FDD9E8CF29DC5149CC674D57D30A764AC0303F5AEEF29F57929081CDB7191BC1AA767A72F7D0F5B36D0C469D95E671E9694A750D725270685CE0A01F8FBE4612F4D34E44E3DF95354DB1BD6F5AEC3832A0017C0D3C10A4F8CB6E529D1633651A6BA179DE2921FAE547A12E275B3BD6AF7DB642E4D8A1C47EB17776EEC4ECD66BD9089B218BA5F8F2F654AEF09F5660324D1779FCAF3E2306D305842214F139F691CD7DCB7E13B6E7A2F222FBA8978435998BDFFEE3783956C40945429D9BE529504798139C09CE2D165D64D884F710285821CE0A1A8A4E29E109C53C40DD4517CAB7F2B8CFDC575795EA8921A21A609945961FE2B3BFD1430057FFE35154179F8F06E2E58055BE680471B9FBCD4E81D0FD2690586CC42EADAD730E7E446BC95FD6567023EB5DBFD5EE8CB6D26D8EB61EC6345F2AB3FDE5FF3ADE43402BACF4BB44277A835D48055C51444652C3598BF0B33A1B39171D7750E9DD7BF0AA011A34EF7A2BE97F7948E16D76483B4EDFCCA6DEFD4145D1D4257000EA0CA63972C2997F95328FF05AFE047FFD0D4C8D884AF673A5737C9A99DA11FA1C446D8DB8EE7AC2D5B389C6305C4269EBDFABE62F9C55578A5F27FD856F332EF8C04CAD67E04FA8E37C19DDA270C2DD70F209DCF90ABA68E1C56E08876E3EEF912C470329B36BE5BCA4E0E9F5372CF857BF6BB45ED45B3FC37660C3D5FC4DD4561F14CF792A8CDCB658A1444A8DDF52994404D542950EA5FBB03DA690124E6DE93B77D489B63C5C84AE595D8A46F0011CF0D6146A371FCDE3AE85B587017B0FA63B9B4A9EFC436F686F1C5262E2447165C4B80B11F499847606C0DD2594CB9100BC3FDEC865C5D4FBF818F3BB95D4A47BBB5A42A27BCBE60A53A054C14F677152D7E83796C03CB0176A86DDDA93E8266B821C9D161E68E8F3C69EF525DD3F82D5F387A3BC3036984860611B64BFBC9958D631F0C23D64DA7BA477CD5875207875EB9D972D310CAD82EECA7AF8D49D6B93E76A4655A56E638AB4E4C8DDB97712DB59FFF21B4080C32C97A630A0EF8F506D5586DF87FBD265EDA8D7BE042935291F6B6A88350AB11AC6F242381B4C1C6262E8E212E2968E45D224FCDC5B47B56ECFB18CBD51F2395F6879660641B49ADA8532F5C99804EA9C28BC7A6E5A29842CF883ECA62691A568A28A27DD32A7024C9356F5EF74BDF2BC67A35EF75AEBD9904698AD44012E318B227A779AC1524F77B3C55A33B9DAC5A5D7EDC4582CC7D32A14E93F722EB611ED8ABFCA3A63DAAA3C0B7BBF2E15FE79861ADBFA131BBC3AECA4EB656B8E5AF362E370323350D071D200E01457A478058A44CDCD2228F55DBCE31B1AE5ACAB1C1FD363A62B88CE43E7FE131879792E07BFC11206AA6AC6D6899BBAF194B87FF519599D85BC37D6AC5B6837E8FF8EF977D4BFD35591C475AD591FDDF22519BC2FE7129762F102C78316B3DB10182FF6679DE01B50D85707B0CC8E8873CAED5036885018E5E69757F000BBBCA985323BD19398EF7540347FFFF88E0A48F2D83EC36D504254018A007D656B855857004EC6C77B4C09B0BD86DAA41A6FE714BD5B960413B9C3F8F34CDFA29032D70F241A68751EF64E6E42D717244B475E59A31D9842948C7178B3D5CDB9AA5C97C4BB15FB68C99A22559E2A90852287DEB10689FF380792251F83220F414BDC88E36C39AC2A0854D39255AFD4B9ABF49AC3171996333FF40E574FF3CDAD3C87F562E43C79CD4AF5DAACBD2F3C15F9651340CF3BC9314F7D1FE606F71FD30190C181B5CE2ECF456A0EE05AD5A05FDA055E5FD6CF3DFE09AB2102FBBF3749D625726D7F161B47C4EA100D39D2DC60701B953E30F5F8740E4097C105E3B9557738B33746206B7F338F55CF433C3EA16C26F6A514AE82995CB89DEA855ED71AB953497874489776C0B9DCB38F453C9C2B2D2FDD0E62A8C0A1277FDDA73C391042D5147FD869CE8C040517CD6F33B0DC963516BE6F19FFDDD311E232D4AB8BE8774BE74011C2C141EB8EF6FE407BE2936A54792314A06C3A253642A9BBAA1AFAF3584941C72B211F583B6EDB54150415CB9DECFF968F30B09DBE6B42E2297D4A6A4B134491AE2147441FA25560F9E8907924C338F4754616ACDAFFF862753F0A80DFD54CA58D4A8ED6D174EC95ED9B8DA6DDB811340E1A3F97C8D1DC3D0828B90C38330C878F6E314607371EA4DDDF7EB72CF09B3E3B42B3DC5CDC13BE80961DE029BA755C52BA9768E64C76C1F68C63EC905CC31618E2C6BD9F5F3226D727827E09053131CC0F13E006A410F1F0533B9EF2FAD6130416F55AFC316B669A9E1D073E7715222B56D7666FD72D0E4DB2EEFAB5DCC4E42EC0F51E376C98937583B723B25EB4EF4DE17BB7EEF4D409353CC794D4E0EA51C1CF55E3566313971EC66B43D0524B0557C3DBA03E86A374B44B814B03A769E0C78785FD540CA32991AA4E92798854B687CB4C3EC1B1E957BCB9E0098CA5415D58E4DC2508C2C093F2AD5217EE603EA4550DF04504B2D5A3BC9EB02490A5D6E3C22CF2A83CA9C4781040E1A75595E66CEE80AF6399137A4B9D08CEDD3AE0D4E444A7BDC4CD1D24F47189687EFE62BC7B6BFB15658A2B9B8FF1CFC5619E360178CFE00A02115257F3E6298F24A37C0B526A5D034C6994D45EB9DF2725011B1DF0BE0BEB09B526D87F377F0A5E7A455F28E4D67CBC26CF84BAF9CF28F9C19F72F087F979F294F028E7192A0BEE4FCE1DD2C8F8B4840BA5EA280E7FF9EE0DE1A9436D5A2C88282811A95A885210F7833AF3AD36DB7AD2D04AA481922AA699737F6B4B03718AB1CB19A4639754564A7BCA292693518D5CE446DED4DE5331CC8540AEDEAC9CB1BC51970EB4385F29AF1F82D4C3E73BEA225E17D7B52DDC58C9CDDCC2C10375CD509E10528D83DB64CC0C0CB1271CFFA95811B24479ED4FCCB414828FAD2B35BBC0B9F1C38083FBD4A281C504FA906D5C5D79EE06BF36874251A0E679587DE68110F74194694D233618618AF13FA16D9A8DDB0D83AC56B3124E6B10A3CA04462D72F4B6683AFB275B0D9A5D7258C5BD6254A08D9EAB6975C75F8C8F90A820D075D3E3C6ED13B23B0B79A8FD221E129ECE0BB8D49A7A2A1149D1CA1A75F6A0F40ABC7B84F793B92B293B07B8BCA3478179F286319C3B8CE168DB6A963EEB76032265A079AF8C91543D5500176B82ECA467F905EC09C359AB262B0198F7F6703952633BA957BF8A8FEE9004F5D6B30C6A64528CBF24C8766E0EF8293A1C8FE4425AE6DA77ED5106E4A82AB4802168935F551E18DC38CB102CDB28FA5EA432AA9310366E6A0261887D3EB57A34E541870946CD7CC712F478B940DCD975DE35AA226FA9C1B861EA1CD1D52BC0B1746109B4AED8844E651A3CD1FEC0542F436DA8FF76FEA5FEF635D1DB1BD1D15FD66779A50C1CE3873511110598C7EE43B538B3B68BA728FE0615C1925FC96F762FD5A9DD141957F72434969FECBC04C7C831947B57F12570449DBE641407BBDBB10DB1AD8FA68559A40BA7B1177D9BC479D5AA1B951083D173398399630C02CBE5BE0D78708EAD625D298BDBD2A8A9C837117016D3A189CE86322C3D08D2833FE78A59B135C2D5E9FC7DBD1EDF0A139F669C7BE64BFA563F6F433B567899E00A486AE5E6380064A307BC0129D0F901C18894D6F8ECDB9ADD6091C19A65EDA5FDA79E17E0CB9C343D8558B1E6C7B6C130EDA1341E9797A8604BB1827C4DEA0BC992D8E0A229FF62CCA37E80853BE68EF30E0F8461A738C6984031D03E68D7AC05EDFDCD56A9DF306202EB476E2FE8921BEFEB43F9EFE9B7502F9A716A6175B7EADCB07DCE026EDE4209744B6E98E632B19C31A410C288B65BBBDFB5882149E65E49D05462AA3E5D83FC1672A645732FD52292A447C3F1CB3113180C6FF2DA688C1A90D1C8CB6554408978128DB9D973C83FA86289C5F0EF2B992FC7FE7ED6FC0EA43C7FB93B5F8D852C6A48B31D6450EB168B36EEE90CB89A4A0D2858FA70AAC22B2FF21AB48A4366975B867E9B3928C188B27F29A9273E964734338EC624E0A2D8E3EC4625D99D85A4E0062792FFDE8D9BFE7DDB2383A6177627E4521FE8569D73297E69B6C4BFF68D92AD5F3EB4BE3B8653772CC253CC575DA30AD5D02B28423F34DC513B64D1031B302EEFDAF3BA80FDC47D383A85D25F7AA9CE87C7CB36BC827852E935BC00038BA1A294B336F11C2AD2A116D7BACA822E120D3B686CA4CDD4D226DC1FD553AEEB54F2F518007177E536E47C891B9EB94462CE996AEB687EA6CAA524BED6531F4F3A3276641EF4FCBB6816D0DB5B8889F6E5A272E4A2D91DDB57041CFD2CEFFC17CFC811A595AEF6E5B34C33F933D5BAD7A251AED27ADF074BD80C0305DABFF7AC1014B106602C589484EDC3BA24F5D76A19F7BD249C1C2C70CE81C1EE338BC386F668EF0B4FC4DF5F763AFE975FD5DDA9EA4681AE36FE150F2FF0DB3F8BDEDF7385138FF29FB1A0AB95E422A12B4C7199B15DBD02FF489A766B8ECCE0706533A8DC19E3C16F8EF7975980F6C164708DECE14BA4BF77AB8D68E4EF8197590A3C9CA59711B93952E5661D24BE8CB18F65ED1615EAAD01E93FFDC32D2444F514CC080DB850DA5DA402DBF8A6A8A7A94096193486AC15023A4506617F5D4C3EDE1CB5DC57DD57989A63B23AFCE746EF916D1079532311DA986FDB0FE964C'
		context:   'F510B36297FB02B4D5B0443B34718E46EFF4E0BA603BD908530BDAB3BC5565A50C2B4864DA1BD4A2BB186C0D7C1AFF563B6F0D27C24B183E758E7E6C9EBDCC42BEC05533C7C9B6FD1CA206797A4F96D277797189982465615F102E9119F045C191E65D12EC77CFACF8A54B28AD774EA31F975DE47E5E281BD241AA9776AFA367CBB3F1C8F2B56AD55DF0E7C03F38A309A7A440BD58117483AF4FC8564C2D9DE0668B605081F5475F55B6F5F3E1D76B9A98F7C4138F0AF32C0373BE3915BF8C52E3C898AAD23C016BB7D0C74C3D78F66D89DD16D88081A9FF3633'
		hashalg:   'none'
		signature: '4E21984D8756144B7D4E419607ED9A3C471912F4584D03F617B782BDE96576AD470606D6B8AD8D4BF016C36653DDAD9509DD1DDEB6A537C497F524D735A8EEC9AC4F582144729FDA2A9625D1C850736CB7590D5791ED933B9A9177E61A4370D8FECC989A0954690F543E77004E854DAB5B11C407CA12200CCBE8B02B643E8BF7B2EA6C2B23AFEC16E9BE0EC928D754E503F2E0350DF92712568D05D4F889A9E4B0C8AACA9D69E71E0AD72D93AA4BAAB5BE23A662DD0B812E81C1E88E9CABD59ABF2C56F8DDCCF1A443A5D83F288E439C4EA18FD26EA60E2B06051CC7A606AD04541DE9A1BB8A49AC6AFDC056E1698CA3C3E4E8C6DE871D4BE04BE8633AE5E5A9D1F62ACE606323BFEF49BF46D28D7DF683ECA490F1E2059419181647124A81D8B327ACE38BBF78918935ED4C38AF2FF41BF3AEC18509E66ECE2200E61E5A177A2ADE2777B8BC526303C8752477BAAFD8825B3288DA3D81072B9F060971AA99C7767E4C2F1BE79A5896DA31BE2A4B7D92233A59548E2D52FBA905951219B82F63FC0EC85C3913CCA3FDB7BCED10DE9E78DB49D71778209D190F03BA3C8785F3DEF4542DD50439DC2B30EB27D4D6CD6254A8BD814BC0DEA53ADEF05F8A137D3E13B3245AD3D0102B814B1395234F85BDD21A8DCD850EE79314E3CD1EBDC9ED0AEE192F81D02B1E75E5F565D0135FB0348E6BB2767F59B439B92FF9F191AE362DE71E106A06CA2EB71455EC1D62C737BADC732C0D70990743282EC7F38CF193A46C2D7823EB4E27EC7C75A5D470B652F534F4154B9D03DB10B829C4A495F581333B3D85D4455C811F496FF4D26ABE1E627F27C350011B53D379297D53DD92D93415763BB7CE1A26879E2BA420B5E42606082709B180B7C0C4B130C5E9408C5FF7B85BB1AD57EA38BC25809CDB6A53AB0C70325117AD5B538CD94FC445144A4A132651D092D3EBB934C9D31079194EAE9874B8719A87AA724D31114C40E6934F7569F7DB681713A6AB4DA36F8F73B76606107F902C2E3A2C86BA39A7B044D08B26DCDEAC1C1CCD1FCEE9409BA6B9C85FDD8899DEE30880245302B1391F94D0D0008CD8A4A6433853C94BF86103DCC54BCB0D8DA3044775624AF761B7D2323C960969065BE4D83ED0CE18310E814823AF76790441DF45E1982C23397361743EA195C4E9FB8FA2EB6000F387A6AB5F69FECF393DC13BB4BDE1922E606BAD7B71FE7E2B0399E19F70AD4BB4E068FF0A7D7741F7A708988B9A2AB7281A068D91C4B10B3963A139A14233B06A87334A1E754AA0BA919C7682419D826085394807C08A7BB3FC8DF119AB0CA59B7CB2DA43FE0556C41175BEB1EDB4ECBD44BE54348030BEAC8151F4BEC2D5C441FCB23B48ABB58C472C7C07680CB6E611DEE2E41D72460BBD179ABFEA50951614D0A5CAC9875BFC7C70602E048A5DE35982F8D24C0443A9FAD5CFC2810784424EE2F500ADC144CAEB39B5402852B83A7F2E859AB261CFE5D0CF6A0DED888290845AF3619B7A52D0903F57F463AE2A06A2328C0E5E27B0F9F1BCDB2D372AE55282AE1D834356EFADD4CA6E11C19B75BEB866F404AFB3E439DAE78B3E65D1DE43A754B2095749840AD8337273BD37E8EB96747C19A864D77554C58BCCB6BC7DFE1E73FB205D9B6C4134AF43F5A28F56CB0D5401DD0245E3E7044A3FCE7562ADA82EE9C11EDA2A4AF7D9B8B8880BD8A5A35D69D83688CE79D38504F16FBAB8A03C61A13F0E9893EFC15EC36F48BDDD444DD3F819020488840EE8B6B3BA1C4C47622FABDCD29D524C58EE1C8C778C286C05FE37E7DDE0BDB80AED0C7932FDABEF4F3109F766AAD4BB95C6EC622E12E001E75031A997F43514F3DC86204978CF0A90813C892B190E27D604816110C062A22DAC6D8E4E78952718C7117AC9C3CC6A29E1984E49F86E919A98809893F02A86D4D45C0CD18E558896E070E8DB117328B27AF6702E539E37884DF92F957C29B479C21B34764035F192161959F0B409827BA01775C05468F8BF9092B07B9293275B865C4B187DC1DEA1728479C126BB9730C34F20131E71F052F4D505C3006F160D441CAB23545AA11C5546D47A0652D93F2ED29A3138C92D951E4CF350F7DA0659996DFBE7D594C41F5A28A9AC75406F3A05CDA5EA49935CF58809919219DBF29EF801C44A7C30F44724C7ABB53B3B2F33C5657E4ADA9D30C0CC324749FC8425EBA88294B3D3C816B962844478C2FCFAE15FBC2F24647011C226065C932E81E60901582F3EA495781FFF509B9329EAA2DC0C158EB0E0FCCC445FB47519FA0AE995F5F5D63C15934CE35B81D8B04C0DB3275CA6248F41E36AC59583FF396A622085DCE07746088B2D3734AED247A93BD931FBAC3509159BB8B3A9A6E95CFE9BE753E200936E3E5B923889A5F08BEB74A8612B18789DD3DE3E99265538E019E65C16094B6E95D585E6671305D9BEBC6F03720BC41A765CF330BF19A15D34CC3625B754B9F66396FCEA2C0A6396686A8CEE533F8FC3773D6641D98F6A80B764902690DBAEE183A11C15BEAB59B35C7FF62DD1AE76EADCC530A4C364FA0CE8B9CCADD3E32C9237EF9FBD690280D0A3B7B7442E56A548F50B797213C26D33257655FF73F17CFF4DD84AD1FCAD2724DFF12050BCCE063F5069F005A41A9F65EF4D86EFBBE3637C51287C157CD9E2F156849A1155445FAEBF5DF3CA2CB66EBA2C2992A713D6A7530568ADF7E2182B9A36BBFBC0F526ADB6C99E38D6D6E09B0857976493B6BA7FE781A0CF8B0FF723EB1341C858A48B700B71E5BF50B758264890B7B539B57FDD65B622437CDE94E4788465E00F502F296B271B6C87451AF1CBC620FB0C1CFD430212245569F385950EC292AFD11E29073E26DD1D3CF4D2A09847FF84ED31910819015CA9801FCFA6EC445FF1BA5CAA8D69318862504C7F29E56A25497A8B1D8FB974834F95C60886FB4A318DF8CF528E0416670B9827DB3511960ACC23BF9B3B0056EAF09B9C16C9B3B10F4816BA32CFE6E89EFDCF617D1557B1921B32256B631C63F5A41F78B5A30941D1DC9F2C451C949654548C8B1D80DBE8DB1CBDF4A922FFAA0DB4BE86586F05F310D5B5C1E9BAA7CD4D630882A0FCB006C6F1857718B830A237E638E25CE6626AFBB0AAEBB0F8A83479B3C2EC89A01E806940F58FE6B346F88334B53DF8A7BCBC4B1C23F12AF67F8DBE2E2857B8FBA2044C09CB6CAE2081F51D8091C7941B4861B7DF9A7D7A986C60E99E0EDFEAF1FFF79277539FCE6B3FE6DDC52ABD0707C5710A4F13740E5D80BA4B5197E256E24A397D5F12118A20FD72E5F6E2C6548334F92C3EF9DBA4A3075A4A7BB6B87B07626C2FF9C3442646C817F34072C996C6CC7488FF257D81B5DF1A2C33815E9F8FCD708D0B67F75735E398CA9924A3D2C0A86A8B6E7C2D738C1B512062AEF9CCA74C4179E6702C684318EF68A7D4FAC2D171EE7E25FCDFCD0F1CFC1F2747037C00E9A20AE42E6DF14440B2A2ED753E0DD67E8E619BFEFA8EC9546F9DEB1CEAA4F26A7DCB9DA79297971A8B264C8B805F1B403B30F5B015BBFA7B38F270C789E928F3F9BB88EDB11D69BA8E712B2775E24D01F9C678EBD301751C597FF1B09FD509E6C8CE8EB4A6EC475A45BD555D568AE5080A503A62469BFC0A8156800FB7A74A1833B10EB86ACD18DF798E57CAC5E75AAF13ADBD468F6F0A4D6537A43366464F9DEB5147EA252FE7EA886CB48E8BBF2AD3829C8824FC26E67CBD8D2CB72468736EBE9EA93A0C654005F808847DE2C293D5F828B0D9A9C73285D7FD7BFD530EC0760B913FC95F65575B3E4D6A81D3C486B3F4D20AAD7CB8053A8B5F8D645746156A1F16930B8052CB4086F170FB010390CAC46A42C6C48C4259524984CAF3D4F5038002B1953709656EE0D6C0E03F7DF45F8BBF726DAD9E03CD9CF6FDF448656F396B5426C6F1A5B8B2B65EBF2D9F3FE8D24B9F061202D576CAE5F32CE7788714C376764CE0CA79B80AD6C486DC2242614A7CA0283D739E0F2697180D503540A44192468846460982278E9586C2CA89A55A3D4F7B04F7E9EE6CD32C33EDA3E54AB6FAC8EC075B8A86033AC02346BBD07E298564AF13F9992E2749088929907592CD51B33E77137164C992B236BF1D73E8BA6FB36DF9F1A40F0299BC306C65C114EAC1578F66416F10A4B94381B34FA2E6CA6A6810B0FD79A22942282138BDF01073B5C9AECFA09E9D2869F0F5B24862E5ED5C4546AF706E3E238D3284D480599A5208FB82408A83E6B5D7D43DABB88781E8B6A6A43B7CD38E493E422558318FF432FC2F35C07BAE05F28CAB587C6A5F5D76D983F50C52D69A566C29170E8C3FB8A09F2FDA97418D0FAFE93D5F2DEEF7B38BDC4B6E95BB851FDB4781524FD9381B981C472DBD1103AA20364486452AC88B439BEEAEB772E0CF01381EEED3ADD1CF6A2063C881E54AAD72CA32E7B650F6C0704051A0D6BC78FD50AA65443E9580D461C7D245002D461F736ABD72625FB9102FBF8C6D727AB68AA9F8755D8C1E346BAD3F274AC917AE1061EEB387CA65EC66136A545C4DA583AC4566F25E9D857EAEB83C9651DBB240F0460C2A2A6C9B2C99F3EAEB3177EE898B8D192E2589C1C5CD309120B20BC8374FE1A438852783B62BF56210A205E096CE91C77B1DF8EE56BDC33E772163A54C9A2E641796FAECDEB8968E6EC45E4BD2EF0FFF5FD7F1EF478D1C8EF0822D38EE5D33D17225AEC4FF62A0444C4E94F73F752556B2FF84EE641D0E5500AE74544B9CF6DA19A3E5FA0C431DCC74F90944A4CB3A418E3EDBC1BA353872DE2BAFE01F8004E31CDFCDF4D18C164397EFA8D623FD9DD007DB14B1CD5A7AEAE18C75332565D0AC6FAF0FC148AD0E13F48EC6D5364F468D3C7160AF37F424A8CA42C8F7A11A67C8A61077C3028B4CEDB1DA8C135000DD822628468A28B04BC41E1A2EDB675C0DB51394725DB29F93E4414CAA7AD28511124A1C82309674D72102EE46A87F16B000A7B7E2BA946BD6115D9F7BE4C8BA85D319D41F84849FDF4DE55D060AE902DB8E217E04950BF5FA96D4FABF33BD121813FC852B0DB897D3F0C8E245D676EB5E41B5DC765BBE9857D439F3C1A4003065C22CBDAE0BD692BF8DA7346FC6D35FAB58C7FD799745A517C208C2397257296E6C00C0A6B8284C0C23565B8C68769E3E8911FC06C4411F4F70E06FA54D4DBDE6DECCC5C5FF6086301ACBAF729FBFC778329DC23E1D1E6D52D86DFA00342906B0A3F7E20348B0D15D8ABC9CAE426BF81B4AF0419B885E9D1F30022477FF1EFE7AF47530C5281C503911279C3CC4BBE3169AEBBF36E56DE426A715DEB913BA2F38542E5DBEEF2621611E131D635BE8D9D1314B3156EC054396656A1628825CCA7528E73BF8F652052F9C9A13CD8DD6BB756B083B4C379C03786FCC79208B34EEEE269AB2501D89EC55F05DF4AA84DA1866E838FB843B92631F32413A3A8E57A0BA12E662D75A37AA1B594BDA9C7EE069587770B4A73A905A153DE93816FDE9BEC16A39DF34E5E679F582369A3179D35820E1FC3162CBE46F8DA5A8EFD2E07B80355FA1BF0AAFD3F12743D0BFF9F03C31360D9587B1178274E257919F42254A87A960296A8B6C1B3F0AF6E57575CC2A627BCC0D34FEE86333CFAE9F38E940E71538E12B43FC8629615ADBDE403A09EB14F67571D573B845330764464BA1875534AE3B960D5BFF9B679D4CB85D644ADE1EC44328D364C05F5AA9AF5C99DB737AFC565EEA90E4FE5DE255E73B48134AA770AB83B90F701088CBD0ABD23E6F327079C10E2549DCC2154C3DC4704545C7F803AB9CEC80274892680B4111E1D72946BDDD42BA3FF3E81744121AEA20D45839E612D466147370384C339B812E684E92520B3A976A348D6F56B3F4FCA8D740D29C7E90431AE085CDCC7EBD997FDC8C80DB2B62B044B11B40855E8A7B1A93F8C8019040BFBC5122E3663896138546F0F23383E66D4A31A5A5E334C7E7C14F3714DE309FE846A75D898CD65D637BB04AB3EB1D3A1F41AD5DAAA745AFE4AF63138B415653F7C25704AB423068758485F3EDD309CA5AF93E5934DE8289ED0B3D65DF81AA4C208CCC8C717359EB8749C11F3EB71BD3A29BC7BD01304BEE2455B0674DA5177A68BFD3FBC431C5964F0A588762A7CB87E26A0F0A13591EE2ADDD246C4F404EEE7D1B9B7E6F3EE9790621B1417A3BAE92C4D32395D8324761A74410F0EE80655B247D9A1D2699FA8AF93F47574420645ADE82A53D4A1E9E618E4EE30A8168DE0DFB29A787C369EE1EE045E790FCB3FC2E53093A0DCA80C34C0F80C29B9AC1C615FBCB5650850B68D625C1832D8204DE34810D58F767C7CB9ED4D307B1C7F87762D71A77942791C48EDB85DF03A430A2F7AB2CBCC081E2841736F765AB7B5F4A91FC94024EFF49A9882FBF312C48868920BF198C2AB9BA6F2385F368393A3725BF7CEEEEFA8D1CD76614D07718F4B97392BB0B6F81335C4EEE6E9A78A445864B775E3C4BBCDFB05E37F15B465CCEDFBCC4F94438191C7889D8E40A1D26E4F39B8E2E2EF0A48EBD5639F20C33F987A3BF9FD20008BDC7E1C03ACAFE8A2A5930977199520E07F06D61DDDD55AFDA1DBA0F5EEBC86D10B3DF85ABD6E89BCEB4C2D45377A690E0B3AF0834FB2F338CD2A21B037B6AAEA6989B93A6E74ED1152FE371EBAE15198D19CA895E324AC495654F604DB99FB7685B5D2F578EA6D086E74695F747C3CFF46C6516E17272573D1A8283E89DAE8A6807588B8409367AEA17E099C5860C573097BDEA7DAA0D0434554C1BB648C9700ADDC5460431CDBFF966CDCB9809F1431CAA9D74E5129B7B7E4C4ACB15865491A44A47393BD58903AC868F2B07FFA176D2BCC902D528E9C209C645C3086DAEDAA6E0CDD14B8D2C402F69CA2E76213DF1B09A6B18C0C004CEE6AEAF5F1BCD4ED5C6BEEFC0D41A9287D0806A56A966EEC116A52CAFCCCFE85685CF3A5CF57F2C959767D252FB4AEE193ACB414D38F5F9E6E40BF0BA9AA16A05092BF3540701F0EBA006BB75913800B3F70BBA276C357AF8D259C788E85687F92E053CA03C6E3B57F87418D2C8A3B9B94978BA4223E988BCA1D27B2DB1569817BA7032AD745BF4D5E1BDF3185400A13ADCC3D1F7B27A2EDAEAA454E0CE5E20620A9209F4089A7FB24E982CCA40B39EA58B42376DDFC59107752E053F9B8AE74E947EB7DA063A9A0378F87441D7EEFC9F2B63B2ACA69BD826E9DA6D71EB4317D812BB51F1D8DB4ED5FB88A2C72510C9D71B2BA03D4CCB7B0D255CD52C5428B1D2088DD53D4C5821B3059B582D35F5D2753A9F6AE275D631790BB8AA010F57C473392CCA753FC77A29C99A4D41FF9513452EF787479C139BA68BB0E5F85855B9CA69C171B131DCC7E62A9347D58CFB4ACFF04E3D656965541965EE667E1877B1D8C7052AF8AEE9FFD8B3C349954CC79BE1896F11C70219A57935228CD2B8BE29BA8FD941A17FB82B8A913990586B4757887A3391B2D4F2421E6F327A5D5D71BBAB42D25D19842CB0832913FAEC6760B6B185EE6E0A00CEBEDA465D4A8A4A673D7F17B363AE00BC28F966D2468EE0CBD98B454B31B759FDFA510BD88663E42B51EDE161D794F4E81B3FA6C5C49456F1106E9F9AD7A7A2DB0DF1B57ED09262252A284369B07DDD8683FC8FDBE70728741A69A16ECE5C486ED980302DD1583C5FFC74D513DC38B594E57C37A3BF35766897361DAC5E6234D391422779A6387685C29BB5E10CC3E30420ADAA8FA6B8B1F89C0102ECCF5E3D3D67393EC8F86D9C2B4BDAEA421FA2E4E4C2815C2E935B128E2178EF99ABC129A311F453BF6ACE019B30A240AC748567D4A7A5CB077C96F0A6349796F2EE967560643056D97CFFD33AFBC13645EFCD3336F7F2ABB2270F4FF466BC08BA5F9089CAC3EAFA7A44C25EB385F50E0E4204DD1AED23C694C48158300DB34B5D40574E4386A25A706FE666C2322203EF5C8B9FD4D6AA746543FCDD3460414953CB471092268DC908CB2F0A74FFA5EF4DE10D3AC4F9804DD465A71794EB70ACB72A6EBFA05ECA6268ABB5D636B2DB00C560D5652981462339AB655DCEC0B57F0F50E612371157FE3CD99799DA2B66D4581F67A053F0D910DD0399A3A1B7D69CBA47B03DA2F184D541C4B800064F4E119D70CD465EA0F66C16E8E1C46F8F9AD982462360C82E30F55E04BF2C368673E57CF82EEDF0F5A1724F5C1CC1DD28FC24CD33CB14FE00AC720E105840DBEA2F005C7B44202BBFA977FB9609F9D5712F7EA7FEE5887E52F2A82D80B6E6A5C7CF7E2DADD4B3A61907F5AC72D315BFA5D4475EA566BC2D9BDD796263E213D5C5B3984D1091093A58DC54F125AD6919CFC147E209BACA59578A252D0B3CFB45B57BCF82492A9B9F29180673E9D6043B9414DC5A859AC7618946E1DCE5DBB6130A7C05C41774FCBF33BEA9275DCD29E4D3A65234A3445A422B8EBDE3B02879F715534D0E48FDC6620BE0EE1AFEE998985086492D68093B788E8B0995410EC3E71862998EBA5A2D12634674BA04B096630173D30BAA8B605DC2C262277A2FAA05E546C4D200AFC0ED48DDF61E13CA1F80772A6FB4415F18DA6ACEE51E582589E62DB7F154DCBC910B72AF5B8F7EFF7AAC89D6CF28857B1950AAA443D2B7FD331606483675B5B073D1E00025EFE60F5AF1FAE5118F1F5F371C28594B7F848A1DE0C6A4F2BC4F62938CC4DCFFD9F1E0AD6099D37CC3945E1C8431A72225512683A28ACF6CFBEC5ED903EB6CA40E1F60839075F4B5286AB5AC6743FD97AF2DC855075FA1E75E06A83EF0DFFEE7AC1663FE2E8960BA2DDA394B7165EBD77D8CA2E062D8FA537F0D0158ACEDB84E602847DFE3062303485AEF32289CDBC56D2B8A840F6D2E78DA9321C6AA00DF075BEB4A0FB4B158BB4D2D70D117441411034763DF291CC70C2E5349C93EF143C7671F364F12E4C7B15DFF73AE533ED4E998041C109C3717EFBD072DC417E6EBCDB094A92015B0FC83192B05CBED51D720F88CF5F8316590A64199C1ADB49219AAC3A7F957786C90435221A87E1163600B2F4DD2543997AF32FAA50A681D1E518FBEEFC22886F24788324E5B48636B7184E5C3F0B1F501FBD797B38671270AFF31A2D1402E35332B2210B15395DFBCEA54FC5AAEB038DED0B6E01D4CC00F3074758AB356CB8760A27AB084F8885E4BFF279B621AE1F10F6E6524972CC9D305A0D7994C9A497A4E7F9BC04D3545C610CEC3E2DCF0ED4FDA25D8AE57EF2E787374CD5C3051041EDD16425CF11108AA3CDD5B387AEE944C12202160B5E681A61DDAC8383E1B90E1C8837FEEFD913D685C63D18D824ED886D5D5599BFBE2B3F96518C0E955C80A7FA2062865B112C0C2F5B68C41FEFF508081D8004B919875951149B6E5792B8B11BB03B5A83A618FFBE1FC9D54EB994E60F1A2A3B9D1B536CC873DF74FF36F0539D0E1FA9D18AD7ABB33EF793E36AB52DDF0DFEC9B4E8172B930CA8A43661F37E635373A7405B417C9742C77C93F3B7547ABA79F9B0F262C0DF75E0CBA5CC4335852097D61CE73BE38AFAE3E62D309151BF553502063255F7A8484F0387A257B5E6E45225063AE4BB8D1B1163A563E0F01849012F4367C88FF8A0DA5582774B8184DF318C6D3658BD309DACFACC55D92ED9B9F7814F0D74BB5850B46698B5A5D3C5A84D6E4DC38535C520E3769C260CF4A7A24BA589042F187239EE486D0CCF396C6A281836641399FFFAE12B322B0AC4CD1E43FD53DBF9239016358274E52A53667D0AA9EE548A4B338EE3BF3BDD81FC256187B1565AE7C942671C3B62AC38E135D819FAC15C913C2D88CD8CF0298BCFECC70867ACD7630C3D88633515A1F9D53AC59706160F42B76B6A8A20866D7DE7405761EE807A1C4718C38986CA654376B7F2063394D6C0C3A3BA5A834E5732E674506ACC561D9FEF05CD25EBBDB82DEEFD9EBBB4578462718C0ADCE26843085986BC14FD4A17F62097D3CCE27219C4AFA5B0C40577362037D95B155966E77A2890E0AD7D0A8CFF41CA1E133F74A66618C750AEAF1C5CF2E38E7781F7AAD226D6466AAB5E7B239670DE6461E7B76B189364BF908EBBCBAE362B072DE83A7FF898D39D003098CC5395A1A79DDB74BBD6DA32D4FD553F938A9F3B2C1556545915F9E95965EDE18CDB6E6E5F669A526EB231A9E0B6DC8194E7BF644378418A9C9A749A5FAB63337FF868F738B73EE6D6B09E90EBFE57552ECEB03F7A9D7EC4AF5CECCBDE840711EED7F20D6B3F3C6429ACEE0D9DC8357D8A29F2744C3AF19197566041F859AF36F0452EE2158BC9B50CFD0CEE03E02112B2A711AA17EEAA2242C07A8DE2FF35CA6F0F4302884C0CDC0A8FD9B6347261DBFB96D18EC90378AC4A5BF34E64E668CF82546191896D4E37A11D16CE7B7D401DC98F609A5AD950EC59F7D5FE0EE13C24D13CD6A9707DC221F8313D97582E0609D8C0715A1F288B6FCF218E24A284AE1D9837AAD3C971A19337DFC11E448FDEC1FD8A35C17D879F394735B9B5534FC69B0FAB6FD3798A72F7AEEC7636563E5A67B09B876369F98A8C0709D37FF2E0EC26F0045615D164D38461888C54DF489935DC0DFF33F3EF93BBEF195BCD8CE240E1FCBA512707DEB93C1CDC36BCE71079D99363BCB6806521343C41465670622E6EC886532D864E576427BC616AA78D932A1C5EF58EA4F971DEDEC07A221847B8AA5DA80D56DD0ECF1430279ACE4D826E73F8BB04D5B0EAF7A1DB188ECA6EA4D2078840530341B54B198343FBEB2D93D2EF5AD3DE247E6E6F4675E4A2BDFEEDDEBB0CC05CAD53675D023A2D6156C1D651019E8410B4F3AD3BFBB666AE5782CD10D55409425874E4A3B04C02807BE74686FDBB30805394AF8553C3DF638988F73F6AB47AD2EB07B1420F3377F88E98B479BA9FD69121186100D7A342C3CC212516491CA1769D247CB6D9B5A7F9D7635107588367ECBC09B12226690ADBE68E9E67416C892949F54C383FB79265DD9DE3EB9E1518CEA482C877F69CAFB989C33EB9330EE6C5C971F221F719E7F643C1F8F38FBA3C17349CEDBC81F3E0FFAE7CF888492B9273C67EACAA0B9BA8A4058298D132198A3162E4E66730A00677CD2A8A55A173B47D0B946D5C962271F8CD385FCA19AFCC94482AFB6F48F18BCEEA8D986DF002ABC5875BDB295963C7BBC3D596879B82EC717EBAA5741598CD2F440F35C12B7B4EE8D3FDF32AAD5F8D8D7DB6788ABB883AB1C43A9ADA445D76C4F64FABDC03BA29F67193841CCB1C935CD95CB9AD6E1BCA90EADD3C149421B63226C066156A883DF1B0BDA8222B7D25BDAB266A30A99C282E50F5501A9B96A66552F09F7E886CF798B70C22E23B59FBB0FB96FCB0C84509D7166A0E88F6B7A0C6425575C33992A75EF647527F1A5FD60D2A7D8BBF80880E58D7F40C1CC51EBF68216E48D446D3BA144B8DE8BB856696DD32DC6D71F70E967729FDD28A4CA6FE7E39A56A558CB754F39DF78061B9BB25798704EDEB6175B942AA37EB5D712B3DCAF41A53BE1A8FFD8B5CB4505505E812840DE9FCE6161DB29EB013FD4CE5FBEC4D43CC60C2910FFC62A02259328B718BC90685A854BDB6E83200BBA1BF01F8E3265DCE91203FAA4FCD4CECF643480A03F1E8B7223D6D4502B5C39345C14940A8ABFC9753244707453BA8B9741D032A93C02B38D790C4F21D4FCB2C6E938772D22247B2F362290BE0DBEF63F6B6DAA76F013F0B300BDAEC4338FEE62050D0743EB65BF529AB514F2217183F8A74D2027DC0928B190BC60F004C287EBB7793F921DCA04F5AE619D4224377C3C6F9721FAD588DCF10DB4F6332E1F39FE0D59C7F5AED7C38C16F0E512944A40C351875959F8AA39FAB33524D80F46D095A55736E0A1F6E5F34FC1B207900439005BCD6F8FB7AE0CC56F0F8509CF9CB7DFDCFD8E510D03BC1CE4CC0A8B748A8B851CA33BF1C81F4B78664EE3FBFC072D3F4F5CF4B1CCA3521E86DA862BC9D33B63E335BA6D3BDD1E8F82681BDFFFBECAB8E83018723D04F6CA5D38D6FF023BE3D513C2D922C421CB7EC2091668D9A1CEFEFAADB7443CA8AC1B9920B251452E1509756A115AC5D04873D00981382F2B8629316BDC7394DAC3E96D01EACAF563F121550E4537F5BDBC19B48B7348C1E55B05577EBE5E81465D939D2A56A4C791C52152B475D6C455E4EDA6AD94A9358D27343EAA9FED7DB7598F40CD2E89FAB5F83A9FCFEA34B0806B83C6243F21CDC4266C8A721EB6DB8FAD4235917906936444339F2B1DB401CA88840BF73FBD9447C7B9C27CAF264992FEBAE76AAB8EE444A0D2816DE56BFA0C1F1EEE7BC067A59C78CFEDD1A4267260458266251D81B1F5AF2BC40F7B6304F7B244E4BB616CF251F62583C56353188E5FD3190C39DBF6F1F657D154B370E462B2F84D9950986BCB8DF6DDD53259853E2BEDE0FA21CAC13499D34C4629E738502C077320C3BDCFD77F6FA7C441EB23AAC11AE7F552C93E7C03E41416630BFEF0C927AD10685DEE67FCCE37662A022F35821200092849539FE32852B61D0CA29C6D207812E2DF98D012938F99D7F72739271778A48C92273535918F6AF10D43DF924BD3CB459634574713D311B9ADBE6A7E6A07BA198EF8A81A8320887ADCCCCE032C3381E4CEB4B09F299D97671D6CF6267D690BF5C213DAFDB1327F0D72A5CEA3E5753D9E32EFCC32B485AFBB2268A63AF9A0F53357EC158D897140C5F41D8750902ECD3794D298C79F5C7FB719844D59762DF413722F43EC3EC0680477395FCFA87D89EC39526C196290581A99022B4F205EB217596FBFA41FC4A513A56FE625D84987A8FED87F3E2DE6F4435CB202DA6DE795EC389C3D2B1EC55B925399336A575FA34273F47F20FE27DFD45AD5D186783343A05BCC7FCD619126FE4A96F8024AC3CFA0927E01C3D131862A4E8052C5813664EC8FE02953C36318B67344879CD26E6B670BF143F0BF2DC9E28F79D32AB38CD95AABE7F0B575E754148EC045A0BA6D3DCD984E2AF38C15452E3A6FF738C3ABC62E49169B1A02421BF3BE39D277B174AAF6C925B84F8E6ECD679DBC827665138522D98F22BBC36D2A07A9CB257BD1179BEBB72CAB348B9EE82E896A6BE179D6FC18B76E2FCE47E2E06B6E56A309E754262F5F78A07F1C705E06D188EDF8B3E965294A720B4E24B86D79DE07F2028EDABC3E5E6C924531B59D2AC2247C9678C7B36F04E6B0DFBB16D4CEC69A7D880B8B74BE739FA153F3EF84C43CEA47E50449B2AF4E2581EE3D3B80CE73A327CCA8D745E8621EFE4255AB3E8D2585F6DE50867D89DBD95E9FD8BBD3B3019C4251B54740ADCC1C0329630F3E69398D8225AED821162B7FC9906F45E5B118A3202B967CC214B18685934763EF6499EED094CF1668B972164F1945DCCD0D5BD51034FCC4E9E14DD2EC8740CC525417905BC47A4735DFA19D91A3F4777EEAFFFEA03D3B25F83F065E4CDC7B7756047B08841984D3EC80E5E813381CD60D2917D667D7C780EC5C1477C5FB23E07E1669FF6E80BDCD981312BEB7A79DDD453E51242339311CCF3BE60B181CCFB35B74F99275322000632230F13CCF13CA795D7BAFF0BB38F1547EEFB64EA5D5702804E0AEC67DEC90DB5432C55C6E4899D291B29729E1CED80924D4A3D2E577E76DBD5C399930A40A15F688F09A08491144C6663852878CA748CF39F224D491B6AC2504BF9E1F7DF99F4EBDCCBFB2B8BBF86779BDCCA14DEF5B0F80539F9E6CFCE7C0CADCB9F0FD73DBF3FDE4B4A8AFB910B043FC9E0394C463A169C96D2074912CDB1517966A07D78D46E73C5F362D6D9A91F22C8D6893EAECBA62676E648AE42022BA287B84766CFB792B82C2A74F59CD22445129A66B6D872AEF7E86BD3E3F48FFEBCD6A6D17B64A4515C3DEAEC3DB875980261780AA06242827FEE4DC85F3225CF54F0DE5369C00C73AB4DB1B7013BFB86671F360F182C3B9BC9132AB5DB46D1150BCC4B8A4175A274272A9E39C1B41AC1D27FC6F70E8F3DC75C9B48A860CAB571A09D26C24C560E89324DCC4A29B12CBD37D06786159213FB8E873951C0055E04738AAF9BCB55498C2FA95A1849B8080D6147BAA91CAD8FF13495C989E93D00EDBE322E37DF74FABD444C8DDA1F18603060FC41401D947C4E48BCA987BB5568EEEF90EF8EC5A0365269BE7059343BA9CA12C218E15ADB51C7FF7B22F7ACC76648C12AD22BF99F3791E8B6DE2861BDAD3B69BC91B4EB4C2CA5418D6B8152F64D418A2ACB6967EDA3C30D4B2FF3829970994750215D33AEBDBC8EA9203B150CEE35279290CDB89D7C8706549D3B3F30CBEF2ACDAA6173CF43E2EECDFFEAED74DEE7809C6FF817C4BB4F40283321149CDA456FC3B52C98AE99ACEA2CE90EAB8389AD0EA7D7DAB649BD5E67D7D405D1FD231027B4F0752A3F72BA5DC3F54610EBB3C116730F06CB0D71A8DE52CF9A793FE8F11C1CC0E234A3139EDB49CBA8398EDB314B80541B590567B7D1A4372B5459A54C6B1324837068AB817DBCE5CA0FEA839EE55C50F77B7B6829EECC020BE85543A163F78BC1E292B921C1D1FE15F8852F9361504754D8084B0EB329E96204AF86ED91B3B9908976752183F9AD594854025D25F761D60ABC8D525F7C406C674EA50214FF975B330FA3615D15094226B2985215194EC6D3B47A921739E73033DD6518A2B967FCFF3527A592157C0EBDE942C97AA130F25D33D0CC3E58DD187ADEDFCEFAC96827D0C2E73E995381327FE891306D18B92884725F0F8636382CFC4E92D785757A0122AF7C9979330E73DEFE2BFCCE939EB785111E8C6F4596D6E8C80CBE481A69517A50C5DEC1F1543ADBDDDE4386DE47FE7ECEA3F9A8DD34ED3D6187BD22A730B655DEC033DE2124B925CF648429C5D532D3187CF6727FE75B0332101BC44CEAE3B18F26784ECEA90AECCD05CBE2D95CA63138BB22987F88D5DEF65FA3B4F6A190A0A7B8AF9046899FFA8659572FCB62AF73DA35620CC6401B4AC7D44DAC8B873936201E98B233D611CAED87474942E8D01764245401BFA25D5ECDA1D5EB4DC42B15C5254BD27BF3A55881162E46D02179E3E861DDD7AC10D2C6494E7E4A490BEB77E0CDBEF3329A4D7DE9F66198DDF01D9EFB194368BA9AEBD6C751B364B7DE499DE6046CB4DE950FB62059051AAC9C4CB22AB26C157CE2C7CEA791C2C26D0D37BFC3171E786DCE0266E3DCDE67EAE3782F5661222AEDB16C269427BE102696104D86937B296F7C2818100AE23FF5C9E3085AA032CCD60C84848F986B05B3702F4C6B3A3A586C9C6C96A1D6BFCACC91357DB9AAAD40DA1AED32AA5F26E665487BF59AF1A23F6EA6968CB05BAA32F1009AA43271EBA9C93DE952A3ED8E33E09ACF59C8790F9E2B6B6862F0CB813E74D847BD1BCC9EF08AF800A3E1EFB8A54A44E84DA0373A6AC33867314D1112B67C2C208C540F57FCFC5F8FD10493135910101E800FA7DC9D3A1C6354003C87F753F74A351A7A19A4979534AAA2093A2D2CAC8896B8D06BD8D7940C4A1DBFB75EA0D1C0C44AD6D9A1095CED8803389A7F0C4CF6B079225D5816F91B1F0FE31B876006CB241F6B3774B1F70498468549CAA3925B4F7C79EC177B007ECA89D62585365344171EEB3C8E57CB4E524B02F0E002A14214802DA35D840A7ACF20EA1082037938106F8A59BF78A5292C3A3067FE84F0BC8ED105F709E3CBC25A89FB6C999B0A912FCB3E29592E4A74D10354BFA63F4AE0B0A4E7FA5BA1234E21F966135CBBAC647C1A1A336AE15303030652BD62268B9B9DEBB0D0326031C0E97D957D21F2F83BE281F2EE3EEF6A892C74B661C35F9FE6F0D88A73A0B038BBADE4C73FE3A1FE691D745A6E09B5DF5447D9FBC3FC4F07336B89E6C65E7467479018BFA655A34010D1A9BFBAF83AAB6CC86F9693BF2963C7799B41BC2EC6D7CA64A621CD06BB5C40F3E87CA9FDC8E1189BFC317E63F6E58B582FFB10BAE2835C0D1972892D476F78E4BAB48B53F6BD5B2B860117719266C1C6405F2EBA2F4F839E027B4EC88249AFC32648B13DA274DF6D86AB4FFA9FF53377406BCD3CEE15961CA76A8BC36FA17FC9CC31F44F34D21D075407B323EF75F4D50604BC99BBAB737ADEBF8463690C3A063A3BEF93745F6D023D3781837084267CC22CDE1FE1A2DDEA2485329D401D6214FA5FF82B11E51A45531AE2E44CCE32126234E58B0518BE17A6FBBE2DB84F25EC259823B7C2978787D66C66DB700A7C20541FD3883113680D123FF52BFDBAAC790C6A67390CF323CE1103CCE0368F96322BB3000434874E8CF87C742355EEE643B39C4DD9D315203AF49C03B561D64702C28863BEDCA5E226336BD63BD337ACC3CE59153CD8F1FD79F42D145CDC2BBAC834F04AA747C4B60146BD4A3B0249B99BFB37B93F7FBE1900FFF2AB02BFC5AFBDAE946933C36AC62FE78B4F1807D587E536205683CE113812841D692972A1387A3BAC9F6820CEFDFE7A14D768D079B5CEA56C092480FF9DD049DB796C1B93384AB56321A18EC99AA6F1A2967D7945F8C1532F9C3A3EF02C774736FA36C8C892FA04EF2660FA0CB90740F1C2F25CC69C3E43E4F5345205D91725631F7659D7263621297CD67557587F88CA64C51A95DBBEAF600455F0FDC87349C7E5A5D82E26AA8F7A4AEAD247838C3A6E72968365FC9632D58496A863E255267DE8FC7FD5AF879350A37A5A7CF5028CDC0696BBF8E5DD0D1D983E6C8556A5C162D72F056BE1299A8F66A9974B978AA4FB69F62636BC905BF55C03B4E3246A01AA1AE091132AD76E7EF501F9468CDA10A6A8C6A9ECD0709502070C51B87D7F47ED27F388C204C9F880EA70DAEB0BEC82B5A5AB74C1CE1190118FA0E060022C61637504E1ADF397BCBF9844A94E97FA4D09AEFD38CBB710E5C86C05719FB02A82593E9C2728D81C04267EB7200CF773C6B4A0FF6BC1E324D366D0732369FF4967C99C3DF28C00CF61336B93A35D191553C826B4A1C6A6804691F95C90E8BA010885843C72909E7D8BC243777186A7C459B1B1B4F8213C4E4703C6853B59F9F123D43A2F81A66A2A8FA00FC49598B464914950C28EA7B3FAC20E76CB5DBFA283C5A67DEADD68D9371405F6596C1A2115F138BF043ED4F374F85EA472B959CC8866BA9D07D627FA874A0EE3525B060FFD777D081EB26A97339536E89B91D2AD862E31486CAF2795EDBF386C2C94CC9018C2AD6BA54E42EA9D9C430C3BA6AC7FF46B98446202FCF112E0B21ED92075148D1F541704A3A45CAC47A9A7DB8FA9C25A210AE808248D680B13071B6FD10EA5FEAD788DAE7C003B77C8638A30E3B0F204F106B2FC44AA2596E29429255D8CEFFB93BEAB8B4F3A21ABFCAD95D8253E33C2ED2EE7FFBEF24BC673C023F4D5174F7BEF267D23A45585B4E19F529502D676A2F5140E4E297AD1902C0EF3F961186CE68A1CD30A2CC4F3EF2F90B2CA2681FD0652FAEB64F5E28CEDF9E2A4B0F1996BDE73979DA7DED743833AF7488C10348430396993736CAC620D7220B02A91CC2E06761442C7B49C9EC206D87AFF67CBA646909B889A997891A90013D25FC03C94CC4DCB8B3C1FB9DC5F334C723B2AF1E32A1DFC19275CA3EF2079FE1EC53C461652BB48422280ADF6953960F5156E01117A4F51323A9E4564D2A51734E22C99BD366BCCFE461A62B8D487C96952A32CBD9B29975E326A9F1BE01D7F8EFD21B5DD3BDC2CF7B4B9CE0833DBE5159B44368B3547E044D066D3299E25A1D1F3F1436DBB793D0AA1DD013FAEE7C352AD192B1941333C1F424486E7144A2AF0FA3352DB436CAB6217EA0B9086489F64A63E095279160A39C95F62D2799975C2F42E84784F4E4EE5D38851AAD3E76B48AD3499AECF071B070EB031714187035D3019C733E326C146F11750B4C12B13575D00602BE6B6F7CC6EE19B680624E3801B537EA56B1FCC20D9061AB84B92869286C102B789399D4B3DFF71EC57BA92DA81400CEF0076DE190D68751247676B69450F21735CD1C10FE373B43B14713238A063A41C392BAD989ACA1535D21D22907AD1187CCE444F4AA55F66271BFB496FF0CBDBC0F17A92A4EC18485B3FE24F4A7808BF4BC9C5DA254D88A7DA15F1CB46815553235F7DCF4C21D170C762E64A758DE2A7C16D27DE9F0FBBD4432DEEC78E40EBD34392F17DDEF18A35CD3EE6B4B64650194210B8FF241AF9F7BA11A985449A2AED7F6F50DD3006E8208AE42DFC8ED9A0173B8946C9DC15844AEB181AF11EBB5125EE15C099F3D52023A9FCF9591CAD15A2F9B4EEC7E19B1C0F55F09CC2B97CECD751BA56E58D75D1E8BDADB48B8FA1B45538D8DDF35ED888190F7BB61BCE36BB5096898BB31C069E8A4DF7D844A70E8E3AD8A02824D8DAB846B4CD7A69CADA8AD8D1F49E844B342E6B267927770F60282D21252A0DAEFF9316E3A0DC730256AFBF73A0CA73371823500862773407623C734FC78FF28F1DA2941C02A25268E831B141826DF96B45089F667BEA25BF05FAF36BE0D550897597DF64B4A0BEA9F6F1888166AF164D573A058A337D7C202E33C1650509CDB42DB7CC344E4257D09CB4ED27B8677B78BBD81C80DCA5C1DF783E47C6B37C35D9AE2FE09102660601D7D2A7DE9042BFCE19E73F0B3BD9B23E6F84737DD8206446F8C96E8946572D643FA4F1216392428A6C95F1B3E013C315071B84E852D903271B9B83A4D582C073C8A0B084F3D0CC7AE74BEF225EF2929371FC28396AB973F5C34381903C25A837C19D3364816B13BE4809A9AC692B9ADFB526486BF176F088CA559E822D6A5F0961B78C78B0FB920AEC1447FD5CD8AC6A809A1333A3ED7A95CEFC9449DD3D7B9E52BD59DB84BF53E25670B1EF0FDB32447B82896F988FD79898FAD3F04A7800A90FDC52B1A3285123830935C12FC3AF7CE7FA85754AA99901DE318BE444AF089D8548289D954FB1819BFCF0039EB2E984CD1F7EA80123BD2336389230E4ECC2F2BDE8CB262DCDBBE20C8D1BE1F4FD248CF7AA89DE01EC75EFCCB45EB337A32B9AAB7D7F70D48CB43DD4DCF1DD95205F4CF4C1FF1D2C0EF9C3B1271B82421D4598AC0936A6F8B22F1E755347CA56ABB4DEB95AC3EB19751645903FBD23F03AC3D22EC14EC13EA86C2930B64FAB330BFE6592C52A12CB68AA5C790B4BDF340E885E94CC6B6545D5F440AA62D3AD676F04C9ABB1DF99CB73EE364551A530B597701917A0ED70E85FB86F4A3EF0C949F7AD3AF7875480A1565E71B85F772E7148ED0011DD287A1428587B52ADD43C33C4380AAC55374FDC36A94F77565078CC081136ED828E6A61B990D92811EE29918441073D1FC273F965699BDA6192C94F1E9462FD2CF22B96A74AA4B8B45C66E5F9F8B296062AAA71699EB00C1DA9D8333CCA58D08A3BC7913E41C97FF00F48F975F737CBEB5E090F4ABC754040B1FF664A474F053D117F7FA71D59C82CB20B23340EFDC57A4351AF117E91A1CC16A4A5BDC64BFBD486964B7D7688A80BEEB2AEED2661136953788FB1AAF531DFAF07D4A21EB3D70E9F9A0877AC9282B25C5CF34E9834A11D62161CC1BE88146F8995A7ACE7A2F83CDAF95AD3B10583602D734074367ECBD5CD5FC25B5F22303F8A0C81773E565261BDC04A8CDC0BAAD96026BACDE7418F6B6EFF7374E95A0E8A83BE8A0E88EF7AC2FB9823A387B7E605E019E8541A4094ADAF5CDB430E60B944C7BA24B901399FDCCF4514FDA7F6EBA922A1810DC47F2065208055B1C63814DE1EAD57A64F3A0F287E3EB1692CA235C10A54690C86AD77C4DE7C22796D8BE2085D0C96FF49634B4E593D20BDA7B8A89EFDBD35B6D5248D3DE298A2F1AE8A184BAC30926A6C97EBAE3FA074881D7F27F07E115380B8FD7491DAA8C2A84F6B6D7D88DEF7AD46781055AB07FA364052AA8EDAB1953338B7C99458E284B846006F8922F7C972EEEC582D3600C45CE0FE7CB90F3F0B68D9C92D865E1209C31000A964C6FAAC5BACAC851F2388D89EACD5A3555738DB7177AEA5B1C63C35849B55164CF223AE5DE01B81974DDB5DF176988434A5B8914343B605AEE0D56899C7D02838C2808A302B840993F24295BAA948E6EB1F4D09C9D013E85894E19DEC8D0F5810AEDD8110A7B801034F45A621559D43774AB27D2576EDF83E2C7937C601803F757972B47E5ED4D9C93F72195C85EF8C2B98D78E0AED590FBCC6B6C6F15A254AEEDC57736C623FF887E7871FBF3817B85A324D2FF7223F788DEB1F13B56B676FACFA03CEC9E62835AECC74E8B28FAD298DE646035A96BAFCAE294EC7B793C5AFC589E4527C31F1A9E7F787E6D2F59751276BB4A1A7EAFC51E93E1A47D1FA0840BCC0EBF675CC4AD11E22F441742927D75FCFAB2A4970C6905621682E78FC017DC3B14B595E2D30A3BFB2C2CE4411BDA084D13907DB102E3B2FAD411010200F4ADCDC03645940B0D98BF8E4AE18B608863FF86B5CD21C4AF05960BEA114F9F873E49EFBD2CD5C4AFFF506B71432EFB0DA221A88968B46157E015BD3BC038A302BC889887123E28884F56535C3C406F9E3466DB871B3FDEB8A9B5B251EE6941E171DA90D420BCB5275A66BFE32C623277331A6E2BD515819459254EEDF1A516B2D1E3E8CC113723E3B56FC2DC0BFB07AC7F5E3940D62A8E075FE8A83504FA56C288F7336FC0D559D1EC8AA5609D15C927C655F805A33B9293A82AC4CB5B84824E42861BDEFF15E0DB5E8F8DAE241C1B480F0F30DF7DD372321ED80071A03C3E853CD8D46F81F078A0F78E0AD3616CE93E75CCB3866CA58788A3476E5D7ABF7398D79033CE7B3989E7DF123C7B3FD3971D87FB51D5FE06E0DE77B8F2BDFECB930C8D0E6D75919DAA0049EF76CD89B0B6B2B6E4005040AF9CEB85315675F41858E1D45ED4890E601D7B2BEFD52C0CA692F3D20E76F8440DAFF0053B226B0FAD4C1EA2772BD9354041B592DC6CBF62B55FDA542D0B50F07E404E7DAC0E697777303FBDE3A34F30FECAE8896AD6745617EFA2093B193757010F5EB720036D82A9A3C7AE9B194B17D767A1650A84C00A7291C91BE3158CDD4877DA8B2CDF4308A1946B2444E4A032CA68B90F88FE1AF78F1BF582E8C557A297E247E3A69ACDC02AFCF8CAC4A3EF8B21E79EAC77D40D2F61F07A8719C4714F28A8BD9996C7B83E078D012F0E0E11F85A415270B752A1606CFD79C526A0FEDEB2E6E1DF56C38A4534E21D6B1AE5DF391690119EAC184109EF644C0E8EBBC9E74B35738D878FECE268800C830B414E9D0C35573971722D0F3358992B9E1F1F273F0C8203D2C846852CFD821519A8D9FDFB73BD851FDFB70B25B270274511A1C0ADCD80589DCC59802A90670250454A6EC5B8B2E2C36E41FEBCAF75DAA0C32660ED5EFED7A1C2FEA55A729765BE43DA55EAC162DB38E8EBBC738C27B1E0D360998D33FBF8038D82C70281ABF38CB4D4F17AC7EB40828D08EC5948A9F47C68963F9E901E9B0DBF109F281F96FF30E80416152E0FA66B286352BD1F0F6F60FC641442CE96650ABFC3A2312F2A2978741997791F9E55D5C22E22905F39EB3DF73333AA358AD79C930A04A8C2CA3633CB50870F1F3D8F49E45D784CF3C0B3FF70A9C5AA51A285F04C90AF001E0A3996698AC7AC1C4CF7AEAFB28CE25AF13BBBF87964FB9A84050C9AEF640853417AA19767824589526179FDFDA6CB0C5E34E1D30D560C1D86F36B0729DE4A508C4812AB9D6EF452A40DEFDA1A2E5B823B2CF81E7450646D3106101C8AAEEE8BCD4F5B3319D6D503A0596177BD2B8CC1AC1A249CE09B6F2423E255ECBAA85C40452DE55759D04B82921374016055FBD2679DF5EC068BC98480C29611997710C77FC66FEF7A3CF9A48E0EA2014D711D86163B768D018F17E815BB794D4467903333367C79ED01B99879218159124FAAFA48A67A30F1EE44FCAFF45BE9D1306D0BD020130E147617DDBC4FA3B6BB97BB91594018A7E05442C30FDFF4F1079405CF09B3C036A03F5D7F14DF937E627BE8BB91D0208E2C8564FD6AB1E097B57A33A354DD270ECF1E2916DC28A1A3CC7A71D812D16CB34641F0CCD0C5FD1F00C694DCA6548138991EF50C459DAC955CF5925362CF91B540047DA991A7B4D58BD93E4EC329FABF0F6B3E3155CFE16CE19DB7EBFE92947BD31CD418C2C06545DCAB8E606FAFE1E0BED4169C71BEFA8FB7EED422A967D0930BFDF80C0812143990172209BE0B3EA734A504CC820DAD4536A7CD4E2324EA0F60765B1D2ACC7BD17EE6DF3490DE273A94211DC26FEC0F5359AAA9756CF2A98E79C69AD3A16E68F41F1FAACF0163723C1FAB76C73B5FA30DAD9B6C0DA2863ACCC80E2609F9529574074684199DAFC21E5221F7147D7AFA1A90991132857E34993CA2BCE3A2B81BD22B2AB251F106C9D2413271DCFEE7C42688673F83F5AB43854F20E365C33E588D5820042419C1655698746D1AA80FE642310799E1CCA2EE7C5ED664E56477390440FB2C63438A79AAE1B8B277FCD0CF204EB5B79B8C3CD73F9136F55999C319FD67519B1DB181867681289466DAED2DCD21CE844AE0E343B2BCDA2D4B29AA8A506F281BBD9C66B736CB8AF20CCDE7C1AA9A12F7F098563F479B64EDA7940AEE4C6FADBF38389E7A66BDA26DBFC1E9B082DCF781F7A4BACB3ABF3EECDA1591902FBD3E6E8DC8A47ACD7D387B604A9CDD84AE921885C131BC2BFE234E8E932251EAF9A3D7BBBE2E4011296B27D37DF10C09DCE68938E929003C9AB299AE56538A14723F1CB8A0546495057718A9E46E9A9A0A9075DE87DD124984B47DA1F284239B0749CB6ED9A9549BE877725C5ED0B1828E1FB6F71312E7959448B7ECD694E40F0E581CBAE3CE08DE11BF13F431413843D770BBAFBA1B18915AA76F6C55929E8D3D06BA9C18889AAC26DAE0CB64FEF0E64393ACF1F61D44005E3694341EE87DCCE8D6A2D4F0C6A05F7AEB09567BF782195574AEA0F93224C5DCD2C5EBB32EFEC36D1DC9B82BCF41429EDADF169B632640B503590828A05F919FDB01C3C934080FE22FC95A18E002186B9ED6E4495DA742E99E70322A1AF7C9D721BA711BEDCA98118CCC738C8BD2DAABBD00D07A8DFA0834C4D92556F41530CFD0359B166132FB07369EAE222EDFF009324E3839043E1F2ED769D4141C8B3329FA53099DBEED068C4D1D1CC3E284A8D125E90F41129457ED5501CA6A804319B5C8C44F22E7772B6F458AFF772DDF59EBC1BB9C59B58AB384861E4BEECBAD0C761E7F9B2D1366CBCA7AAF3F2C277E3586665AF04CDA9C8F4FDF45BA0E1EF9EBC620483417494539EE7EB9F578CA58B067C0C49A51DC79003F66C4EDD10C6E8E756AAD36F874069EE8E0F7690E954F4274C48D3735760ABF217C1F3A1216132153D0389B63981F7C4B06951001933D441CF6C4B1E73FF219445DC86578D4E903C0EA3E2E1315A2122921237BFCB2447A528CC28AAED027DBF67535FF1E71424AEE1BFFC3AD28999D075649645299F4B1FF29B89363661DE496D82EF0D5F90EBD6212512340B3F37A568767FBF270F0CA7B620B9DC49A2DC8DB92C0471EEA6B0BE302C9C0474147C3F807CE4389AB25D997A66A6B8AB8C95EBFC16B1FAB6932A5E7053DB19EB0CAB8911D571F392953C49F8F264811660FC84B17F830356DE9CCC1D02C5C55C49A4A4A086558265599D6F4BB9C646133B2289B95CE7E891DC6065BCB356519B9197E382553EDA2DAA396533380B56FE97367CDB73AEC54016FB7FD38EBAEF3076270DE73B915691CF2B1C33035B2C60BB9A7134E39E7EA3FC6386FEF87D9F42668CB2E7E93317F71183F09A51A59A9B7E5793183AAE942829702E287A434409354ED2F3AAE470F6687D4AC7AE7ECBF3FE929595F937512EA635791D1DE34B99E72B2D9CBAEB3812273DBC5BC6A30F80368EFDCA38ACBBAA3D5CF79CACC515E2D7196E2EF3B6BF8B7657298453A0A54443E6F90E2E540791F904E1144E2CB54680837E32694D9FE617E764B4A280DF576959342FDBAE891625AC3F3FF25ACEDFDAC6DA2670EBC4D005122D6C6665E7834B5380BBF57CF2107E2AADAFC7F97C0B16BB36184DD955285D9E35D8FD7D00920AC1F4E59903F232D7EFCB7427DA532215F291400E32467ED008C63C2B6C7D5A92A93F4D48A127CB66C064CFD90F6682085D50A961E265319CE90662DFA99FAE77957EE468B8F60F79C0D1FCF3AA451C0ED5DEFF653EDA365188DB72611F3B60B20D1B887591D186098CF6C84CD324FD403C31B2A539958761A3528A7383B21E51E18E19BCB46C4F7062FB531E1D710966B1F25193D3AA1953BF08A576EB1E68054422DBE6F'
	}, */
	SigGenTest{
		tcid:      1
		kind:      'SLH-DSA-SHA2-128f'
		iface:     'external'
		sk:        'D5213BA4BB6470F1B9EDA88CBC94E6277A58A951EF7F2B81461DBAC41B5A6B83FA495FB834DEFEA7CC96A81309479135A67029E90668C5A58B96E60111491F3D'
		addrnd:    ''
		message:   '3F'
		context:   ''
		hashalg:   'none'
		signature: 'BD40E6D66893F38D5C5FAD99E4885329925BB207D49E62BCB9B1C4685154A8B32E58B70C7AED0E28507F31B49EC7ED6ED6DCB8DB2DA90FE938994D75C80E6712F2421C22DEF8AF88906B768333E7EBF6DDF7B84DC01F06731DD640CF93F57927BB56F9DA9D4B2ABE60C81D863A20F8E5C5CCE74326D6181D01B74E3CD7F794A98B4ED7A791A1B77C561A6E7AE64E4E17481DE4CE7E26065D90AE21C965FEBA3302102D7564E3B7414E1AA62271E9B4DFB42C57C44726AF6FE7F3BDD486D7D578B4B4BA8EBC1F5D7243F94D2D2D4CB55B7F95C3020E05A6CCBE12CBDFFD6466B5B34369FA56839A0E05AF5C6613E4A229895CF5A834880A2C3937CC759F3673567F39FF2B8A0613EEE33963B06D200181F3FE69B507F2172E459B989A8819C7EBBA3AAF31F9D589DC0123012B787B60DCE3DA8A76D1A3476EF08FB8ACB72F6C1F7C8B6929642822EAA13965D6C1F3C58B600CF029758C41E26E0EDB6FD5F2EB13EB91D95ED3AB976E5C6DFE1C80879B8BE68DBFB9F8E2E60D822D88DCAD48EF2EF89F5486FCE1506002E7A7AD8F0E58374E3F82B6E72CF0CD04B86BBB9F261BEA70C785521BA607B8A2DE642C6EB84F691307618C60AD713F7B10857D28613A6418DD1297544671091668F5E8EF5ED296DF37CC6E45B36F261A66B4AD8BF55C63298A6FD79B9A128D44DF4818E613B783DD8D8116DFAB297F520163A15F35A4B96105D7A695C723F11E38964C05F5840AD333FBCF1862B2BFD0433D645F411E73C6434480E7C55EBD1B4E1B786A7A333B8FFC5E77CB303A3D093FA0D18DD223FD3CC352EDD11F95200A2D6791011B40EF6CCEAC57842961CDF74DCC5CE09B219A615B08A9BB92E2F001B7E5FD87D092BE800DFFA75D1D10AD80E543A7809384C8C857780D66B9A7A9A7B15F72C1AEC5EE6F8CAF7D6B128DFD34E26AC6F5267052557E2AF504BB5E8110F28B8CB3268900D37E5E53A2642FF7AD1EC4B690A99BD62A3883537E3D77F80B09D27DB2A28DA659A3B100E3B65088E837826FA707E8E39149056C3BB13D957486964351D88CE1BCB69968C85690C959992AF98609AF5ED34A681FD32F8D1A5E219D38D4CC228182697C9389B2E9B5059B8AC4A280DFE3D6838D879830643CFF92CA02A1C9EB1643516A31C55E0E8D0F9CBF16D01FC0B8CA214259DED8CAEA43A013A645F9CE5300520066CD2AC04BAF8D49AE7694D40BB60AAD324569690218FE19DFA58EF73D62A831501AA25F7EFB5FC9C8150955FE6524DE636CE526B100A29E6E48EE047F33BA6C0BA5ABD5E5720945796A57FC389CAA1755A339F6C584B13D6971833C9E865398C8BF486A5F99EDC9E5D69A04BA1118A3A9140CD52A951D283242B5583282DD5CA1AFC867C14947F68F8D3D91105AC4AA565650430BA9334FA8A8C5B76BAB24D1BE6BBAC8A478B89EF8E9E8B33BF38CFDFFA1D07F984036BB5D9A71031A67050BF451468D1622AD99EBFD71B7ADF09D1C5599C347A8778776E7D9DF5495728FA6E8C6A18FFD7DD6CF2CA7BBCC84B12EE03D9AC24F2EE35F4925161D41F61EC3D51D9A96A1CD67C84E7350DE302CCBBE3BD56EB1B1682FD60DC5EFC1AF97A9A8AF08F088E9B561221111CF29E63A3E7715C84BB0B9756FD8D8A92CAA2EF658E268DE024A54B9B6EBDC681AB04415F5656315B35055160DB4083D184893E8D4C870B803394BAB5E38F5C390FAFECD22B052EE4461A624587F6EBE70B90A840540F009715B0AAE502D2811BB7E345FF2F4F779AE981287BFB96B9A73B999D7778FC47718D47907F60B273C37DD1E7ADF6FAE38F6BC5F392927F18E742CFCBE81C0A4C8C75403361F1BA7F867DD94F4D22AD03C38D554BD9E4DE497ED63C156BA9086F4C8B4D087529EDCC0295A93AFB5373BF46BD04B2E5EA5863C850C3283B3E7524BD5E2ED5937742062EC144E829BFFCB9DAB3F9C4C5DDFE8AFE51BB58BA2D0C8C32393AE9F49764ECF7BBBEE807B98EF8FA9B18A88731B5388C717F321BD4761A74606226C5C9E3E203BF47B1724DA6AA13FF7267B99CE68523050523FC4B8A42FDFAD0F4A0EC0340BB6C1A58B4DB63C03589632485496407B90169AE9F7C7B287E0841B6CE570942FA518CCD80A355F64FD5F739BCC31BAD3C618B591F0CDE79614388B538EFCCE119B0884A850FBA18BA41F39F08E84D8E6B38D7760A39DCCCAF4A031EAE014C6D6188FE0333D166719D275BB56056EA4B8203673F08BB5C44C57B209AB57C17475E22E55B06453998F919557582959376745FA1E348E9DA508CF2E96FB4FEB4B903B36385251B34F319D9ABE258E0B8318A7C9D45647F99CD4A317A9CF017ED9B341C1FD501426BB6C04E12CFB5220AE2A1DFC02DFA2BE4AC859F837EAA1FF14D99D86A26FBE346F869BA7B662EE5B69FD1B8D16FE352BC5720F402A009C649DAE7DDF6CEF84DD2251D5F97C91ACEA5326DBFDF4CE695B5C5908B43EAA79EC1670D75665991AEF8979747976173A5875C912FFF4EE76EB2FFAC233B77FD330B6F888CF0393FA381328BD9936A977DE7240772876BF15A3009ADFD2AB9870B49E79201AB912D57FC237F1D83B63D8EB1EF7EC1055B6A4D2755BCE09D9F2BED40D36033360CB9375A3A5EF8BA045A816914D3489DF7B6B2A2FDB5FADC6B3E1A9CF4063D06B43D7ED75A8C78674CE7858FEC0ECAB11E1A041FF986A904BD84968F299419DF5F960C2736E75718008F9DFCECDF20EA3C9A79190AB27033989A40D3B97D89FF662E63CC0B639E77FD3E983239D8E59F0585B12C803E1BD3A5865D1D4D3F022ADB4DEEE488F2D2C08F1997D8601D702CD9E27984E171A6364C6887E8A625A23EF4988FBC6888A2A49C17CB596E4C415BF2CE9EA4741BD00E65AE90B8C53866CA49F20E575A31F011D22ED8DE7A41F71BD9BB9F7CE42E0A5705C3498415C0CE462558366B00DADD9DA6F17C666D46695B250E651965E814EC70D78C507E4EDB965678C1F80CDA6C7CFD720FC133582F03F848849B261892696765F327DBF653CC7C88FA9ECE9CC172B2E91FFE90CAACC876BC26E44B2A4FEF46A4E2BAD72A55D268E4E99B95D13A196FE6ABF7DEECE54C7677813EB04AF9601B323FD27D90D8701EBF06E539796E68D320BDD2A8638029C6612C519CC44D1AA2BABE31DDAB3A83714C805B98731329CD1FADA30E7E690B949E2E7417975BD83D8130DE44D186A90D0F435C78FC4EB6A02ED891FD1C67BB4052A6339CD75AD525D8F84B4CEB33900F7D1214C44B1EB05C224CC9569FD58CA77EA9193E591E658058E50555C63D98F8528467F134468426304D9771346AEDD3D072059103000906D1843B19B23490070DD6A9F5C6185C34ED9CB73CBFF1599662727CE40795CBB8FC3BB669F670FEC731A226AE12B08FA4F6C23B3C3B2366490CC023C4BE2766168E776F1C186DDE099DAAC158D2CC085577271F7965545F2FF9EB02C670E5CF5625722A140E96291246E941E0B9D0F94C05E66C9EAC61A1E6D5265B9491D6E0FE13C3DAF44BD6AE2C3868E262767AD21106831FC99101E3A8F47127FCBE648A6CFDF841686B27706456E9BDAAE54E5689EC2FB6274749C955AC62892B62AF27ECA451EA199D565891C8C11E36F24B13A74A46D5194272FEB4689F598D2BE372BCA45E177B80D7C352AB598AC0EE6F72C9531074F98860AF8E7D0F49258F50414525715262D689B13164EEC4B8A0419B5E6E1C831249375F6BAB546102CA90333B15A24E543A2579B074EF40E9237150561405804FCA0095D5C4D8D6456DF31DD847F517C8FBEEA4CA8EA88CCE339A4C7A565C43674BD55C58521E4E50E837A76C34CC1F625AEA9D4AE909BADA0C37B5E47CB26562BE2E37402D2210A82CA8E397CB2B88453A2F0FE779E7C6A74FA32B80A99352790B6D871470BA75506F8E6CF0D7F9DF4716D86FBA40D2F2FB7C3C6ECCE2B534B4F693BD5A6DD7E1DA3A1B1209A17FEB7E9830E67BEC26F277921D048F32B9ABED990AB2A7ADA21374D1BD64D3EBC5333F437492D12D5E89798AA7B83E6467BF69E221705CB06CE8B2C96AE7F8D0B41AF3DB1F183ABC5151C02C3CFED01F58266E3C2E67A232DD2D11F8573B670A974CE7D9C8F6FAB7D70C7437A0A0EA38F094A0908F5162E3C63C6FE09701D4AB6EBEDDDF8CB52D8EFF8C174A051A841FC36DF127501B2DA18F087B98B0F80DEE70CB7670066219289E9CA9C1A9EFFDBE14DE19D20850D98149CFF50314B91891097FAA023D699009BCE636E401610E24667AC3D5B41ADADD82872FB0874BC42593134086538DB3CBCA27BF7B8CED845B9FB7A005E813E38971F36BB793E96CBF65CE3E4BB2B20FAE2DFBF63B84962B7D7960BDCAEEC39FFE5587586C5A4E080C4E3C9A370BA4822637524925A4AD8565771E1EF566641773410C6EDBECFEA9382E9B19EAEB05DF8851220DC24B4211D5AD427B8B4824ADE2BF31983B2B426D7E872C205A0132C6D413B53CF4B975CE36749A75994589C34ACC9A87B8B147DC886CC30E02355C84579C64C1D9A466A44BDB6BABED60D143CD89FC9AAAB0B400154E4FB1AE0915A720C8B5BB56875EE54F44ACB9BDB8D447D64A407956FCE1C700CB86F014F398A34466C4F8F8D9DB8B8EEB16762A02B314A05799E7DCE5C1738EAFC729BF655E351E3CD6F061CA4CF25E98FFB486B6DCCAD82FAE13896B7DFF055C58B2B7643D40257EC1FA091C654FBE16338A02276AF20EAB9A21993DDECDBFF5C7F00EE9FC7EE9E5AA5C50C43F657C7E65B4D865B1822EA0CFA3010F310CA66174EB341C82E22D797A252C6A8DE77452E8CC6117673B10041E8165ACA650B5A6DBCBE29601BC570C13C7D8DD57679ED3F9D459F4BF0A29BDD476FAC13CC4CFCD9A3C65B63F57A93DB350BDABCF697F069DD909B4808176E265BB268FB9BC4200B83BC7B18D43DAC8997BF4834A14C4107F3C9E597F77AD3313E670159D94ADBC46DA1F2B69642B7FA8E1EBFFC228A222F951BE0ADF61422878E4939EA32B83242692A140D80DF11D95734E69B952FF7C6716E0B360BE4D0BC3D675E0CFB721681911BBF5AD8040A24901159B1D805CE023E731CCDE39E2B38F096578C9A974AC0CE9A28D923515C1FD369CDA5F3FA35E7358EFDB91A0771F3DAA64E685F5E24BC819C93486B2871FE59A0A2749A15BCFE36C4AB4AC2ED4803015FAF8BD4C309EE883D4F58131F778FBB608F07C3FB62E588CC47902B6A0C646676640AB0EE1B342537E9376CE5A328A052F8F91D66A4AB9A12263BB3184367731930B4789490BF4594EF7A01636BB2775A33E8FD6BF252DFBB4FAA2C310B1130FC0443BECA6E04CF2CEC263B42B26FC0529C5BBDD2643D44F57A392273866626DAC471CA18F115B4346E850D98268BB992FA11733E5F01D2A5753C2E3163F4BAB64F9A19E719D07BDFC51176A327851A7320DA9F9A1A11E57B6D374E26C131BC9D94630F9CE23EA9AD40466A0C6823E0AB5F3282B109B2485B211AD9F62A79E842B963D3E9399EBDFC60DFF8B12266920886CA26F214048FDBCE5282E652DD4C7F0C48A9F8B9935512A89182F81777BE6D4B5FBAFE895DBB4319D32EFC6069A02B87C4CDFEF1955FD3D808442C966E13631A269D206C5CEFE96C2E67FC8E1229FC99EBDCA89AA803C94052973D560F50EE33E74574B5B208A237E2A83DEF9E15356054251A5804577C024153B42C589249B630A9B49C3825B5B41925388A4976F1217C169291FD65A10A275BFE81BAE5C1CDF39539049B38DA2F4FB87E7824F2A983DA6A4FE9B4FE5B26649D6BBF0A81BA862C90648BF8D8376CFAA81BB9F97B080BBE5C6E899B8C9743144DDC8CFB705588DC63741355DC691C7F58D73C9D9E528784BB43E59D669CD7540BB0D8C33EA9C879DE8CB549EB0454172409F95B0F97E3069328AEDCC2518461D870B4C9B7D8606405E46609A8AC9B9A53A0C57B02D4FB15EC8C6B6FC31369522E2BA2FF870606598F5BC5877BDA4198F0618262265BCBE6506BEBCFB463E92AEA4CE08660AB55A3008385AE75FA4746EA8DDE051B9900AAB1F5015F0EDAC6F6C4AAB0FEA3741512BC254E9E2D07C1EB010C88378FEAE0988EF4202EEA1238ADA11135D085225F2C8B976E473AFB04EE2801DA342B7FE35FEA3966F79C4D167D5AEE5E885C5418DD14A91A06032916FE34EDC40BE2AD9F5505BE80404F62810EBDF8A7C96FF7DFBFCCDC32FBE13A03F2D074848495AB0D766D5B35BDD5A841B566A901D371BCDA153F52A146AC59897F5F1BA49D7233BC43452252646C15612F5F27741A97D6C72E892E58DAAE7F6B81E8E3286746211F530A2C302CB4AEEA63242BD6800313ED6F5EF007971FA3DA5810BA9E5F6C98B1637C846AC89E22112A998DA631364715FDA957DB016EF26A6E4535A2B3F3FCBED6468D65806619F42FB514C7BBBF7F08C1A15266253815367014E9B08EEA76641566073879C11B9C6A760544F852CC35705956BD40BEE059AAA1E6AD6E1AF24F26F48CFBB37416A10B146CE0DA60AF7148ED9E8171D6ABD085312AB72CD03979D7477552018A2DCE6164C3BB358A1B7687D613A82ADC25D74D39E72F5BBF136C8C7A82CB3A7A1E0559E50ECDFF699C8CE3D6E9005E03E035075C04AD101CC85C5EE7EDE82880DF1764350A49DDA44C6FBA1E6DEBD083A48F7E94238470AFE01AF6CE430E05822114F24EA0B85541D93F99C414C1385BBFA4745B4EA0B3FB45A94B3D7FD0D6A5FE05C2F32616059621A636ADBE9E8BFFCD4139B0D5A0B6698EAECB449D60E531B8BCFD634D4832499B36A2216F1FEB7B939CA80AE87672E4A7468889F17C88F529E9EA74E1CF1504E81A2D516B0F2ED4794A5E21FD4B9CF5B039FC5FB0F8F77C55CD927BF157ABBA24274D8214A1A825C2F3C8D252FB2B765AAA0A3BEFF0DA54CBC829529E19B02347B8F91BB92813756C8413B6DD145C0146B0C77CC9D01C6FCEEE99A84C28E3A77A14B0B75B56AE8A648F8091DDC917C4EEAF777CC4FAA4F3F9D117CB0F0DB6BB300E913737A7620D1BCEFDA18DE324BAA0F1867EEDE9F7002D495C8AE27F2EF4164782A04BDF46AE627817330DF16094F3E29EC837AE2AF472B867FD9D7F6AC4BF058868AC15D0B7F0D84A639B4A71F9E04E4B4E84982D8E07D0C2C54B78E711E0710F6DD52DB394E3B311A38B64AE960D72E2A655E798C16E7F8D48559B9454DBBA942721350ED975EA4CCAD19C0E422EB9E269117EA62FF7FAD2F8D75561271661B2788E2B2DC1202C5E306BF777107B53A9D65C7800DCED403946E98631211DA326F5B213CEAB5093C5D2E4E2054D50DDE8AC2E42425BD3ABAAA88F4CBDA59B926684FF8D0F588BEE61822CD88360F8EE2A8E55BADF99D6CE950F3FEF895CD8DA4941848B468E4A3C388500D808CF32673417271AF4C6044C4DCA635198D4B924B15BCFC80CEA2B97939575D0D4B6A36F3F8EECEC9BAE05B2A61165E99714A7136C802AF01380DB9E8E504A96BFD015B7E01867193E26B6BAB469B47552C3F4D46DB07340F51B5FA9435AB04113595D786A3409E7E891AD64F154C8A98463FB7AF7BEE76A185B9B7C0EEBF5C7C1F6D5EEE1EC5DDC66F041569FE35B1E343264096F8C567D90F68E21F5B4143D1436A1577169CF42BA5D7516BBFBB74C96112BD80FAD78568711780022F2C679B90E39B97AE28714288890D75F4EAE850C606A38608A23968A7A09A1766F596AFD753AAB473EC5BCDE5BEEE72CA957FFFE47035036E6234C69771D472FF664A3952F9947737B4A119646D646914701EDF2E0DDC4F929F02AC36B1677E49743BF1D715520966696872A9ADE1A5115B9C4A6BFCB40F70BB88AD2ADE2FFC4E5CCA5EC3DBE84EA5AFEA71626AD0BD8BF493006E9782FF67BA6574AFFEC666D368C8E75D9B28BA769246ED84B2D2D1F3240F4906255175837309BBCA09CC6A37AAD50696EF57E6405C1B79F72B866912C17C0C79DC22819BD4389FC43505D78E5DADB0870AE822B4422B034197248E347F8A7B23ED9BA7E86A8C8F3B8C7FC1FCA347BB2295D799FCF603C4A34272D8118421D50FE596EFDF6231B3BF8D5CC4FCB91D4AA5A7719710B6B1AA41FE7FB810FC398A87CA557ED09D56F72D2E413E558A7EE4443A1D48DE20D8F11598BB000FD0CE59F1864BF06B28D154DC2368F57549EC37241DAF9DD776623B79B9C02B81C31C187B65CF29381BD9B9A6963C30ACA466A8DC355CCD024F16626C84D1619BC617FEF6EDC8FA322DD7E0666C9FA6543847AB8222C4325F24232375B7CFAF667E16F76295295472CA29A74391C3484B024A22DBB02D4A12997C106DF0B1EE051017F8D7D20FFE8DEA674CB700CB6056436B5D80F5E25C9EDFA20973DE2C27BDBB1BF858DDF98B33A34EF25080F628400383310439E4E9C8D1782310C23832B63A1545E8D645B65ABA9D88091371808116631BEE7DBD8DA64F7090CDFEB0CBB402E152B3B65773064AB4349CF6C88E426BB6AA51C8E1A80096258767E6B67878C69C5FE0E2C3573ED65D28FC99BEC39132E2ED1BEF3D212E7C36B8F2738F723F4CE7A6D482185F569B2D69F64E719C73CC07F2DE9C8AC3F198C928EEDF178559CBC19C01B925291A2227E5277A00DC4D0FA68A2836E9D0EDE7BBB6B70FCD8216C5CDFFBEC4118A8BDB117EE10833B44D64AD1C672201B593ACACFCCC4AA2C599DCEBC44F37D4328BD82DB4D8D6B452854C08BAAAF96AAE79AAD1198206C803E7196E95A2F2A9E443D3AD1D71F18658DE5470E0C2ECFC4264D34EDEFACD6DBF02CB27127623E38653D3102F3FEDF61817EB2FBD5F134485CF4CEDCBFADB96F4AECC890BE352A3E318C8D57BD1A7618F0DF5952F5CEE62E95731AC62BA1D0BC1B5C6D4589904C5CA2235EFB2D6C2681A6E7C1D276907DFCC7C876352AF7CBB3DC347016AD7C6B8E7ACE5F6FC975C8EEE2F71B037539B2919A0C3F505FB7E91C2F7F70EDDFAE0B86CFB6AF6965061C4D5B2F5C6AB570E891890FA92B056A052B0A1E7EBE18123D14F64BDCC9579FEC83AA214AC5B85F416338BCFF924D247E99ABE3293D8DF2C10A80DD1D354974B2D0972E4EE19793C6F079BB7A7BB913691DE12FF5F147868047632B1186D5C069F9CBA7ED09BD98CFF31DA8698D7ECEEB7A12FCA381619BBFE33A1A0DE2C8B14AAAE85FF17133373C365B198DFE65B3D4326B6CA8188C35F1FF4EE5CEF215C3AD3744BB53A56B1FE8AF8B408C2CEF1F32A6BF35BC4DD4B391787C2E27B51D7E49EAD873A3E4E393008BA1F7CA45DC27B89D8F39F8AD12149FFEACE5D518BE2D6D74F93A36F82C69936D048798DE5E11456D198E617D6596BFD26686451205246889429D67B68BD28D8DDF3CEA2DD5169FB58B64446171A5CE7E8FD79846CC92B69DD03B04468D57FE75CF4B0792093CC1F7AC7BE6E4708EE636DB61F0D0BEAAF4ACA0129D09C4DA407C7BFCF1C7FF1EACEB064F0D8D541E97BA8500FDA615751DD2320F211940EA2060AF8E1DE9661B107C239DB9E866555F85B1DA367940B45792CAF93523D8375C7F9AC2EC5246B3567AD3A3E30668B0A64A29DC828A8F7F7D0F68603757661D3E30A3195344D1AB9126B0CF0DE7E9CE603E75915B45CD1E1A1178EBBD96EEC5FCD2B21B4208B32F3A55B2C89D5DABBC1B62FF40D0004D34CF8E49A2BC2D7650BDDA3523C1EDB98B404BA87CF2D55A52922E6837E5510B782E28BE3AD4B67737CB9656F0F15CE3B189BB1CDB4B6DA5B3927E289B464742D295F04520C7DE50C3B710472B5DA75F58B272C609EB918D8F564382DAC244F2BF9F48CCFF77205114F72900E6BE86AFD590044E8F26DF81CCE3A57A4A7A6FAA427411078BF40289B4E76A18AF73CB9CC44DE82512D74E3804E0599AA2660F949FC52A832AF6EFFEC09A9FBE9CA05A418337CC237D6B5DF9DBE12FE1867A8E41FA87513AC0C29FF675C0A3DE70A86D50E6FF8CAD5BEDEFF0083D2C74326E250AADCA2CE44A3BD4F0A410BD17385E6CA87D3ED1685FD4FFD92AE8FE47512D2B7226A0CA2CE859CA4D0920BD48EE0E629DB896A5869B193F4D4C02D5BC1DEA3B8B1A6A182FDAAF8BC165016BF0B2A95571CD84EA116BB333C37AF7F915ED5C02A307B3D6CDABB71CE3314AF36B19ED69986785DA64AA1D2419F2A4D569C69181047DD14A9C3E112B7AB7BFA8C5BF4B14DDB0226D1E318B0E3319430067D5E4419E051B0B9AA6B126DF7F7685F7A947802656E7D41B87FD62DC509E2DC36D7253D5652B33DB837F6932C116580CF2EAEC35FDDF000C49344CE1FE3ABE380AC6FBF174E9C57DB14498EF251C3C69DFCEF50F29CFBE783F28444882C998454A751E9D2F256252F6B1C12C5B177E64B3D297D3B78A2363B3D2B6E1AA4C5408CB414FECAAA1228BB014384D753A2154DC0B13CD1181AC4C78EEA7819375916EAC65FBD67C83FEAF1397BED4F7489C4CDFCBCF838E3FB72581A832B6B7F1494DF2F56535E7AD488DFB6677730162C34A130ECBD7D70B725CAF6F17060528E24C90A161D15DE7DF2EF10EBB82B0CC830DFC1E0E28C9412288529EA94C9C4D3E60FE2FBED0CEFF2AB6C09DF3CAEFD5D1936A9E99C9BDE73A94E84B80BFF870FE6FF8A79EB03ADF7DC0571E666FC6D645FCBDC5E3D3A00AE3E24B82D18F45BED70CDF38C3965914CF564184AD3994369F436990A44CEB40ABDE9737D160911EF4EDCBCF24107CC6E47047A49ACA096F84CB2BE19B97E388F5028E821B4951AF61AC4FA8A4E1DDFBA6A53C189BEED5493684ED4BEA514AD69A65FD4F29E3E4DA216319773E5EB1D0B42FC7C7DB488266AD4CF48C7C3CF4A229FB1F31DFEF70E0984D933CE90E8567C92313213FB725EF5DE07CFAD01366B2645E9059FB0DF2F31508015D6EAD9E964E94CC93A6FDE5315AD5D6607C3D8C2DA588D06E0FDE261C4A98E9BF9FD6AF3422E607C4D2A3027D56ED8B0795F93852A8B9EAFFF06FADD041A7AF1DA0376D3F19ADB5C81FD513AA9BA6AB822AD4D625D2946EE17B0CD6DB8F4E01D6B98BB535078C72E3783F55BAD3662858F686E8724B78E5EAF7CF7EBF5AC6B35F4E9F59C7FD514F7AFCC10A783594EB1979F37D6684DD323FE90851C4FE394E79A4369281F1C9912A54CF5A6EA56A9F951F9996FCF2E08DD2F3866772CBD6E9CCAE5ADD5D6D180352E254E4695A307C71F65C45443F0DBC59C2F46647E02A29FA767C646A7C432A9EADC144D488B5BC40761B1B4EB10E09147656C3A3C7D3E549F668FCDD41E61002C15797901FC7D6A7E2F6C1A6BA3326AFF9B185E0CA3C312F5661D90BE182FE46BC759405776E08950EB5C3CD327EC52B01C3AEB7B54B9BA3FBB7D4C66B303E8D272D06C3E8483DD928830D604837BE6E8D4B9628DB505F9E233CF8A4639457681E0E9210AB311241F54AEC6A0BAC8177A6298BA585460E035B65812E98CD314845BB172CB645AEBD6BF058510DBAA67098E074E2B2840B3AD835CB58687502BE064B590354433BF3B31A71C706349A4B1A5CF11C9CA8AB67AFC33C69666BE07AC9DB04F4C214CBEC76C24B015DA97301D6D247319F9E5BD48361DE1F460F02274C7D6CB8D9FBA8147BA3750000FD04E353DF79206C47BF8148175C97B068480A40A9CC5EF2F46702FA25B0159F5E666A6605735CE0CB7E96236C84A6D571A381E5C78997FA8EB0CC9CA632295772F699C6744D9BCF5611DB9ECC71BC62790E8F427ACAA966DDEA6A565F0AFC2E05531F5B437E577E642EB390145385511B22901710BBC1C754B24CC60CBC594B316ADC8DD247DE2B9429F383045E0B4A3AF730AD0D34C09E9BC408E6ABC4318D516C9930CAAC7D3544278AC174DC22C089E5DB40AF8FE33EAC9417064BE0AFB8BA64BCFCB15D12B12F29B8A605BD26DACB023591E2C439DA8058B0D8770C3AA1734404D4944515227FE63C3B1566CEF9ED9319B09115F2C5E3A2A2D24F3B39BE9EC6791B0DD736ABA33ACB1A56D64E5215918EE86E66B8FEA89B9F0EC366AE139416811DEAA92BDAD797BB8A81C9B90913ECD79A794EABE510FFBC6441AB4A6450EE3ED1E7E90FEA4043AE945D36F2F1B83EE1FEF6AB31682DCB2755893C0A27D05DB584EAB64680A8BB3D38F8EBB4EEE6FB85DB0597C419622B4F7F0A657ECDECBECB56590C6B6F20BB6D4622C851820DC3E772444066E89F939F5B3CC9E0BCE4ABC3B1550E15416F5718319C279129E8A8734D557949EEE8608ADD8233EA8F48D30FE3B1252EF8CDD90AA548CE25BCD13DB505E2EE5E4866FD6A66F3A95895D487431B0EE268E5C43B0B79E605C80D08DC6D8EC6902CC56A5A78ADC002B16655939AD60353781617FAC8056B79A50E80DE88A52AEC69E22FFE28B823DF1FE2CBE9963CBA9C70385D1D0670B2823364B6B9E633A2210DBDB7516E60F22898DEF3F24545B3D6B9C2C73F2C086F5DC68FE73BA5DE35D4D9E3BF973B9F411EBE65608EEC1727C2A1CD90ADE60DE5C4F35E7934D767AC187AD8C54F92F9E3BAEE15528F52E3EF8125056157CDCA91ADCCC71BC6BC77ED3487FB176924D28348638BF02455B137B66A50F6C8F3872996FA6CAC3C3E83A5416E87D4389D28F4A41B5AEA51F182E4A4D9FA444858D169451E2C2CFBC4E0EDC733EE05207F758A319218F5D140097334A705844DC63D61AEE52003E5A674F7563A7DEAC6B54F93F2C7340C4AFEEF2232143FEE8CB0BD3C218D682B1219C13262665BC85D015AE65771EE6FAA39B4F58F0E7AFB1C90B9FD42C8C6C864ED1F9E8AFE0D08AB7611DC6231B6A2BEC4DF3F3EA10D9C099A6E4F6D41570E3BC17DA7897B78F7FE7E7112A1658972D31D5BA31C91A8B0ABAC7E5443F284C0D76F0A8713633E7E4DD2F4D936C98B479035228372FF093282FE0C22608185F18439907DD2B7647ABB1EDFBEDFE19E5C544723C9D4B49F5D1EFD65E4F51EDDB06322D378B73718F2A63B9ECA920A120F8709DC7A3F52F5351BC004B6CA08230D3FED7BDC366EF841A0E2C788D7B803056BD8B0BA92395A2AA9C446665BA77659A3C3A29DFE8C77FD77CA1BB79A0EB5E861ED0AB23A3C2E9DA14E6668EF03A18295805C3F3402CAB06403707423B6B4FB13523DF22D57A1E5595BFBDE7155B3EDB890B41F2DE52099E3B779D5EDFFB99980BE963DD13E71426EC98580FF1AFB85E50A55C1A6786F583820EF4D3771DFBD24E306DBDB5358829F5D8C9510EB9B0361F246EDD78EC3DFED505D51AF3787BBCD96EC8617BD672AAFB63939016543661B0518A0A1DDF8BF0C121B07749767E9E1CD70880846CD1002C0BA06D6BD0D8468823985F6ACB51362A766EA40F8267B0BB79572B5D9F2BE12873908F2927E08391A5270271ED25396A93BFA994EB3FA55D779FF42546FBA72349157577E67A87A97D4020E455E252505E3EA2D33EE56ED74AC7224CAA24A65DC803AC33CB419EB7415A9846F4DE767A134247AEB27062ECCB01DB51CC8633F661F9F1F1C66A0242D0D017DE5C46951C604B6E7CE2EE4EB7E28C4E9DA71E87137AE236AAE702406003604C0945FBC49A68F55D36DC5F5AE9C5FF8C617BE64F592E23CC5A878DA7EA68C823BDA36755F9B3677045B1FE1D33CCBE7FAE98309F0688DB55951F1334216F4BD68898537354A1D315766EF063C9F19DCA292002F58EFC135D47F81C385C61EE36DDFF51C4722F3B94A7B6F520466F55C327A82E424C340A0ADC426C8474B3D32E257491B8CB0BBDB4247EFE7928370AA7706CEF0AD5EB2D049C6EB69259B45C46E737E96D292EAF346D5045DAA4B81220D748DFE302FCB2A8018A8A1F77E32F6E8CFAA33D952CED8F090E928977F08BF1961D07FD8968C9A7114C5F2F180616BC0176858B1AA2C78DAB2AABCEC9E2C6E0D0E6785579BECB9FFFDA409E9E9719B1D961F25FC7F6791356883DA6B302C44C4E2BB9A7C6EBD72CCBB61669B476E82B5E1C27B319A83248E669B62967D3C94D18E0945EF47355F86B0EFC0242B526686F4230FA3DE5856232BC2D74BA2C7E43A684DB82B8D38BF5D76F4204D3B18C1EF928B160CD139E66EA9F1A619A2871B2E3D7D62A21C30156CDFC2631024A42946E655E5EC7CB31202AF99BE088065F3920E511831E483C75EEC489DEF905B82B6ADE1E8D15D31DCA4E492EFE66EB2ACDE2AF033950AC525B0B2D5429E47BE106DAB0D69000D9903ED88CE61DA1358821D6C560EBBAEE5DCB21063A68C94903D1A58367830D1696C5B915DD95007BB0E97C5D200997AB525190E59AB466B477B2FB940C00E0475459A984F351A14CBB610EF96BE2C92A03749D5C8D697E3391D4F83F5D2F0CFB0CB6734FBC0776A2B3AA5DE85F011B8EF100A2FF2EFDFFCD39691BA637B49BF7E3EE5585D0946292B5556773DAB67075B77C334D40DE0D278FF2671084CFE0A1E27E5517A00CD572EC57FBECA8B4CA4788AF28476D661B1AEF5A8827F015B36B1A6C5C21A23748F9156D2DD6530607FA8AD491FE2FCF9C55C49764B4425F6AD99338FE7F66C65F1259FC9734F7B1F37A92F4115F76C98DF5F7DF73F98CA99C9622E47A91BDEF7CA74EE76BFCF472D8CA9761027004AA297275AA8DE2DA73A31A29E104CDE47E75BDB0B9742CF647AAA4A7343E156571D5002FBE95CCF20FFB9993E38134542F19060A969B9A9FD20CDC01975DB4DA89B9357396521ED0BFECAB974C4A8114030317B10C41B3F12BC6CEEB3EC28746D6891497E0BA38E3077C1C77786153C616BEC2C9E23F00918D904DDCF1E7EE510713528224E87E6A1D3BC001266AD1899AC695CAF7489AF83EA4829593ADE85B7615EE220EC6EEDF7ECF17B5A1AC620FAAF18BA36FE8B62EB31AD9168C104CB56ECC1B2239CE108E403815E47034639EC602AB94630B97995226C166C36052D6B9DBE8955B1F5F7E0B0AF03AB798EE0478E6CD45544503ED86A980AF2EAFF29D8478FB84F26BB230D295B05F089046252331680206E8DB7D6FAD6BC6580862E492193DA4111DD7E8D8ACBD4DFBC6ED2A29418A414DDE900220F9E511B632C9FFCE26B74D02366426EFDE60E49582DE4F9676A660AC778F8D4FD8E616A25433249890264D7E17356E781559E7424EEF88B8835B83B43A0C64DF1CE9A8B7F59D26C96EFBBCE496DE95EB623A021EC17C2A7215A4419F0938DB66D50CA545CDF0AF1A3E5435AD5DBD38CC9F5F60A8F63B5876D90F627312271806C3556F5C910A9F1D75946ACF0912973106695F9DEB91CDAD986FFBE934B0181C6A29BEED3A3B58EBF112BDB94FCD0F7F95D80B7D76E460D64183D5BB91282F892E0070381F95AEB4F54E49B6BD4ED9D67838EB5F24FE1DF043A67B7ED2324EE84268CEECE84F474696548BDB082AEFE3AA0217B9B173E8CC737742584579628000C6FEA7DA90EA1B8A42DD042BE882C7B9CDF46176B6D25F2E4C68CF9FAC5C057E0358E7F919E04347F4C0334C649E21886E599A8C397C0463FC946E907F6E3B84B86094D53A26A22F7A5758ADF1F8841C56327285A1F7EF63CDBA363F3CEC79A6119F1AC8AF46E1206819EB22F7622376ADB62E02601225BE0F05A43664316CFEF8850D53BF670A4171EA3A5F203D5FAD5958E4BF2F047FBC62414337207926F6606098ECEB2DE480A97DB39D1521C10B421C63B4332668EFF48E9C49DDE0A3BF435857BD58B5E5BE3BD0CDDEC75016EDB7DEE2AFFB43AE55CD0359C6E2E41FA6E473B4A31BF8C060518363A1633A334292EC40BFE76887F470FE2032D8EC83DBC7F11FBBDF71D24C23ABAF737D1E068C79643CDC876B768BCA0CFF22988ADEC340D83778B2C72E0C606D7F145343A30E90BBA6002CD3C281BECF18507EF408BA1C231E7FE3BA3205C061813D75CE3062F7268D77570544763CFB5146E648720EFC6FF1ECE9DBC731D09BFEFC8950435DEEEAFE6A3253C40B8A504617F6F1786A3A9DB2E3DF2A62A7FE7F429172CC1A71A3B05FF7AC2FEA89D89F0365823896190F6F7772A485DFDBB9AB7975766874A5D36669FC3A6CE70880729BF959D1455C228E0D9D92C9C24BFFE4361346E46CF617DC746D5685D8D4ECDE45C0B6B93F1CB4E6263BD0B62646C0C3952E5B22821418196D6D79A93C79C1211825C3EB8CFAFFAFD708512C3AC280B9454CC95B0381E48550A0B82FB675B092DABEE19B5B04052BB9F45448B490EFED211A375FAE6E3E090874E0D318B1E23ED6F9527D54DF1D393768B8B990CDCA88368F132D03136EC2A314BA50EE0ABF0ACB381F7896F1974897DE2A17026A72B11CDB4B9F51CCC9D93EF82739EBD6E5C9992CB6A816B244ABB48747C73F7051C90A72EF136BF582F7E3533537F1230B2552D83A63924C7406F5E26507EB54E53729078828E130FA2A83EDAC54C25A49389960B87818EC79160E06B177B869E3D074B621A095F3553B5422AF1D11E1785A0D048B9D13272E9175754B57389517920721C144D636EE1959E9883E06D1D051644E183C48EC06801A776E12E54715AE4B7543E04C71D7644DB759F08204BA5A7DDFFDC20F4C47213B2AF0953544F23B82FE4C7DC24BC0E98065209A9325677B58E6B2EB77FB6D92427B7DD99225C3CE4F000875FF55733AC2D268F9C472405122F66D141260A570D3BA488A7D2CF79080DC1B685AFAD0E4419C8CFE7162823904F2535E6DE0546231E58E368123AAAF934E2DD560BEDAD34935B6B318EE52A7E9B084D11095357E08E525E47903275664836E920E31947634433A0F8C5BA9ECE2825EA4752A0191F2F691ACD942397982E68C6247B9FA1A989C2C897A65CFEB0A0B1827B63B35CA7A1517085B0EBD3C83DD272EAE3C33193FE3D3AB4D1E07F0447128BC1F9D545367E639405ABCBB902D72623D4C6158BEF4304F62B43772DC646CD9EF9CFBB7F221778BD5FCAC281D2FB86A3DC4AAAB1B2629DD8268A9117D2D7911DAB67535D417FA4F457123A3FF7C19AEB95A051214EE18C87239B3B82922F86349E4210A59B0BF96A089604F0A3E7B3C9668185FCB94889366B9B36AAAF934AB305F4F8B69AF39026BD79A57B492D55C1D1FF8C41A3918076FE81B90E3731254596F64D03187917FFF425B142F9DBBFA6C2AE6D6D6C343BEF7214978F7FBC8D112A8595CBFD8040688F304D82130D8F65D396192239EAEB2BEA497A75F889B0999B2DDA23F56B013C7D23893987CFDCCA37E781416F63F8BBEB28C0820CFAE1255141ACAF17E29F314BFD6005E29A322A46D614D2C279BFB688456D028E084991553D2D607368C54ECC14DEC228A1C682C5A450958D28349DA5D024CB9DCF0B41DE0114B10CCC4367857672C86C13059D9318113222D3B4FEB0E2D4A95FA850A3918E0B4E17C81442210140C09F569D3A855C67170C3CBE96F363D9A08FC573DA8D93883F4F270DA5911B8A5C2B6B9DD677CE6E7744DD0E91BB62226B4F8558D06A244969C4694F5AEE49C202C28D33C737DE079713A55EB4FE792F8718F13879129B8BA14EF85F1A97A6AC7A5BB105CCB6E8612B036F3B5F6BD0FB298818F76D90204734A422BE53854DC53F951868E3326A0777BEC4A77594633026BE0BF46FBBE046FDF438968157E95A3B9454BE725AEA44DCB35651882F44AA821E7CB512B2D4D14FD3919A288035EB139501747085527616A8F40F0FAA6B0A4837943E2138BC682A14804666D069633CAB49111A1888BC9AF37E95515F4734B18D119DB48D07431E2D9D49F66FDEACDE44B55407DBE2AA06FE1993BA41ADEF17E1F04812BACB43B7483B932603FC9D8E3325407227232BAC2D4882B68EF5D7882DA8120DBF2C65234DA4685C1005351E6B0993BE819699BF4EFB7B72BDF23C44106B207DEE25BE89F05E4161C828925E39B55DF20E95FC9A23E9F8F6FE6EB98548E3A74C5B09EF86B638D6DB6D8B0183D71595F23687A5FDAEF27E6EAFE109AEC416A7C50DBDFC9E08F1E2033E18CEFFFE3EE18E6AE71D0975983D50BCC9072FA049591C7AB653EC9198C5B4F2724ACC278BA80D26644CAEF85688ABE8D031F0A44A844668BA1F919FB86C577A406F4F4DF3953287238256E3C106D59F701313F79D9E44259A22B002325FA8B7A3105478C373D10236A1FBB1C703D01826585CB925F69450C825B91E0E7D815DE41F411426F18D873DF80052244C6BA4DCED9641FA0F5A8E93A9C84A1BEB6AE11092470CEED4CDB77504CBCFB422FDE56EAEBACB599BD73977FBD7DC1EEF692DC6510BCC0D673484E35E13871E2A8EA47F171C1DAC808276AF1597EAFF6F8ECD89DA10A3E2A3FC6BC2774B3780AD3EDFEB0B952028CB198B18EF2B209FA98B4CCCFCF559BFFBC2E473776D1AD3CA98C40590823E851E114774A565EC690C293211DD869F1AC50B8F4349D9422CF013BD89FF8373D1F39C3F97A6367B116135E16BCB8B57948DB100F441D05762DF0040CD52F4E8C78BBE39E69B502CB99946C4F03A16D1130CB08F378725C10A38461BAF72AD1C708061CC192081886E87CB5A52B532B3E5A0800D02C0F4ECE2BCF300438F96DDEAC6BCAD50A7E3C07682B3772849BF7752A81D36C8AEF83714265210EB6309277C6B866249A8B28232795E05AC93289E65054E096663619CFB208BD742A8CD043BC3BF699D86448589C680493ABA11FF063038C84D6FDAE68B8847C6B35A05C054EEECC4619D7B2EFABDC05C604DA9CD07CAF10C39F05DB6E536BEBF1133F9023751120BDB1720E72771DD68D8000F0424C3B8A047A806433662FF54074391F230239706F27DC7010EB95D1A378121276EFB4F80A33617439F55A1D5A63803AC05C3D60DF8B79EA7C36EDDC12772780CB3637AFFCF391CD154C670590296455B68BB9B90877D25FE6A1C46AD5EEC7B7DA2DABBF5DFB85D7DA34E679CA2C08B60C2F00996CBEA3059D4DDA01880A99BC41CB1A340DA8CE3D5F8C4EAEA6696AD4ADEBE8CA748E082D5A718221CDBBD2058A8EE944A0AACC0855DD06C97A79A293BCE45998100D8F605C023EF62208230511EA3A8F7DCCCE835822E687DDCA1853693A82F3D1C3F090EBDE6E5384C680384ADC2122BD517AAD6D385E637219188D9F11E47EEB948F16AF692DD809B1CDD7B20ACCCAA20E6D1F4FD5692A2D09494231705DF5AA1AD5BF2BA19845FAD91A3096ED81E7ED859D31A7BA329EC5ADCD1F58F89AB2D0963D67569670545668A579FE44B9E1621ADD5C9378B7AFC2F96716FA19220EC93A88C2D551DFC15EBB8BCB4B2B2D491DFDA4E0EBDEA9055A76548E90DA126550F147D8D81BCD265BF10D6DCC0F0893C87ABBDFD545C5B7B6ED2EAB2483650892E011D40EA39202AE8975457ABE4B30E889C8D4D2291DE341976075A3D589A089058B57A661DA35D4E0ADBBF4A98C9107A6ECB8EB85EB71C8581ADEB27B170AA519CD3DD2950B33955EAD57FF7DD08761135EF6DD12251BF92B8EECC59F97ECE985174FF6A81B0F850F927DC8D09DD3FF982C902D1A09D3FEB3622E92EAE2BB9D2ABBB7924EDA2A6E980033D2509D8634917308B6438EAFBCE06F48536DB1D25CB015C65D895F7967E3333ACA04C431031C2E952853BCF922D2A2795E18E2993CE6B123BA928404713D82964FC814B6AD6999FD313F225CC6C404D72FF29522A8FBF5801A3478F99D0648336124179BF91D5D8013D881AB41BD2988EA0E49B2E972A2DEC6DCEE4F3A5553C388E447235F71F2D157C84BCC0AA4EDCDA855057C24BDB1E144C7F6BBAFF79A3DE357E3AF462664A81F9BC503022573F9BCA397AEADD23D6D8F3D312481523F42ADE0BD764B3DA1D6A8BAA21EAFF1CA37228F600F0111A6E885107284B373ED361FC80CF0E6DADE3DC9561331559316FE4E23F7E54E0547131ABD886CE17A8B1B42A8EEA20F6F834D523CE45A069F86A2DB50C279DEBF2965F880BA0D84DBF07A2F66BA4CAB6381C01E4F9AD49587BDF4DEF24590C213D4A6554352FD5815BF24D11A735EEC099FC5EA7828C33C5890BCCA196011E2AC5B65A35F2FE4C361E520DC326A8CD49DA285D634242FB78B2C1CD634DB0F104E510D82852D5494F20CF91B1D890116A535D7E5A31850F648E80FDEDA46E830645321A169DFE34575F1071F6692984DB528FDB9745E5D165E9903E3A548B75EE8F1CA74B63A757EB21A8C33C99491AE0851EF9AE859C53A22B7F182F1DD01AF9645FBB7D0AB06DC14AD717731DFBFEF754004ADA3C8DDD2B15B19C83466D51A2277915D3E112811A36CF1BE8105F592C6EB7D86CA9FC56F0700E13CC3C6B125E8BC7E0DD5552AD4CA81531D7187391BAB9D9EB2B1D4BA7DCA702ACCEC91247C981BC28AF71325C1F1621FB7ED3E786FE2947DFDF56FDA8062DD81A9FB49F386575A1BCA60CC35A8AEC0B27A4CF3E8A57631D03E75F581B8028CBD830D2EFD90B2DE408644B01355D07A20FC7128FE08EFB41B3D1174715C485B5416599E0BEE7B96BEC9828E5D1A1A37D10F2387229E92C9C94B9D3AFAACF86531802B72BE362B9CFA378D752E55A6500602EE54B6B925D8EBAC97B5C032C0EE302911EBFD1F0C9F96485B0D4C20606DD1E5D909EB898124CBE9F9F59CCB7C0186337AFCAB364174E9D85BCE1A12E9D0B8608412E9C1E36268002B0F6EFA78A9DB3535CE4C67C4658B87F3DF348581BB21ED73C90CAE966457A527B0A699E8A762C8ECA17F75981D1B92C6F5D907E856921DFE5ED59370D8DB709E58FDA1C84CAB859D2BB8987B9F6BFA2B9678AF879A1D54EEF7DC7250C3DC4D6FE4C16ADE97D1CAD6C4F2AFEB8A2010F29A3FB8D488A8FD3EF6E07B6994BD6BE0281AC64A690B12594C854892BFACE17941E4F8FB53CE7B7803AFF0BC027E7CA6C43544057F33EB84071F53B5C707F8CFB8FC7ECFDA740B8241F9AC8DB2C2D8665B85E0578940FBDE90A07188C24F848A970EFE1B29E40B69C2C5AB11A2FDEA9DD0E9D234E14647E2ACC55A4732D1C15B7CB014C20EAEE4A46A242D22E5645E0E1A71CB2DA037C69177A450870A9B7641DCCDB2543A1A82FC77522D4FC2B58755A621D43D6AB676A70C9063632A8BD02C1BC404808123E883EF06D5C929C8AC71DB21B3D60DE974349CF5CFCFDE47CDD035DAC85DFB71EA504E77B249120E3F0EB199CC360863710350E076F12D7C2EB7A374DCEE91B159A8C658867D3AF3FD91EB71C9A137F81E54C58D94ABA2978440F7435BABA3DDC081CA9BE505BF96862C6680C487F24DE49A964C91AFB7ED42725E4C103C2626FA85B529856064A9479732A1D7766F5E88D6664B656A3BE1AA674429E0613CCFBBD5AE61D2F4F8A442FA678F58CFD57A187531A47017915767C997E7141986C1486E14035128F7DA92DE3E00508F1D78F3D73FCCD31068C5F518BA3EFB0CBBB8BA3CFF43935930DB7E73185CAFBED82A80D4BCD8D49E1D2B33BD4E0C1CE7E9EFDFEA0A4C8EB10DD94BD51B690BCFCB017ECE3AC73D0097AB44656B0307FE59B7EE626891D1064C29BB779600AC190192DBF462B57E8920366ED252BFF0FF406A6F72D5DA29716CDDC81D3318F0D8E440DD4AD4A5895DA7C8F8C46FF651603AD2B016761663DD7EA0B758A3DC019F3136F9C0385BDEB7875CA5DCA95C74B13F5FBE9CDF4C373142A5B7D348F4AA58FE830F84CAC5CB1A08F9A2E2BF9C1FB2C624D27CADA4599AA5FC861CE933116BEF79B2B73A1CF030F21B04C1BE2CBE2F0AFAEB6D172F255BBC1F04A511B9D00ED74A66DA84B0F1345A4C874ECA97088EC76E717F2E83F50E7E8710F72356B9AD9EC53613C4FE6052CAA6D998DCF470D957E50B94DDC8985FBA9B5D81665CAA6FD5027F0496B2095502442909C4032A477E4CA0CDACBE3EAB381562ADDD43CDD61D4228CF613397EEB81B8202A2B2CDD5C1C5A4645BBC5BD1CCD7386CD382E86D7CD3228F6687145BDA56D3FE2F3E538B9887B5EAEACBC33EC79F6EE5CB92617C4BD7C8A1D8A709EA64C05D9387A3C4D95F36F4042DC87DBBCD9910E45C391C6F4D13A23C47932634C784CE7A96F631015AEFC4C9C4FA8CD06B6442D51A612D270E5BD322E8CDF4B7CC7AE4482AEA324CF3AFC10963C78077627761E3421D14620D95C8953FCAC8E485EE05FA653955DFF93C6160F242108F83065E0BF1367847DF7D0D7300FD5A397D99C37AEFF6905894E19FCDF9F6C75AA07171F0215028D265E5337A37630EEAB770A61D5F9E8F8D5E8E3B46211215B9E246096730E57D75A1357F97ACC365EA96DDEB75FE7EB6B39393565CFB417FCCF5223D0F981AB48466DC16759B02458F242DD0DDD4A357048AF6A5E82F7C173324E84C1952A078AC85BDA36C05E713D340DF854716D7618F712879B573FB8B68FD2E47F8846EBB1C3D66069DF055D92F9CFFD6345197D7A9BD0F7B76BE7CE5021512550BE79F3B2D2878F6B884643BAFF933EDF1CF8CC4897725BFE4A9C84F721964CEB1D56F40BAFD9A0EAE122EA0076622A4464907C4C384D5310F276077C3B77277B9F6ECA541FDC5F1682C57751BA38C14DFFB4D28959FD25391AF503264708B385C311CF538733B18363A7292DE553A9BBC41DADED8B7B4D0A213EC6A748EACC37CBDDBB91F4A67B025591E16845708260344B8B95E01FB93019D3DFFF742BE6D6CB642C870964F0D47DC3A794B38C635C25A413DE6E14CC5B4C5F6A19A1EDB9889F57FA8BA3B4025AD2658007C5BE0E11CCD43DE6AF9F750473E7178FFD9C2A8C212B2AF3CB2AECB2605ABD981853EE019FAE50748B504B40F8BE10339D97F9CD901FAA583E7446CD60657E9ADA31739799D2E07223001F2EB7D96CCD4FEA537FC8630D7874CCD1E4DFC1B763249D452DC959A4B953380F8A481CB2151DABB2973ABD3AF676096E4B1DAE64700F04DF7E80F765E927ECAB9745C7214EF55D65BD6B1D31A00ACDF3F81404BF32244E99ED5554208AD9C6952568C7ED96762123E0FA0E5E02C82C6CF5463891D4DBADBC80A8311F77F07BEC4DBCB71F875B373A8F46E4DA0DAD38622D7CDF2842D621CC1B8A6CFAA85C5427E52B4B3145151E203DAD62399CB266343C396D6FD913661DBD599862572A53C1C8BCF412BE600649C991157AE3288933819F70D6497E10670EC18EE8E07E58E5CE3E686DD5602AAFEFADE329E44F0938C7961E95DAFAA7935891251A62F32F0237E920A23B4A458B7F7932F144FC0CFFCA01F1B5345CB9F9552FBE69FC87E083302C6F0E153693A0715D0BDA2BBBCCF0A48D2C5D586F72B171938B880DDDBBB13DD970D6B475DD0CB8640D27F823BA44272149A7B70E8509B6B574D7213E9EE767AFB9C2242D6B70D0728F3FCEB1EFEA46BB1A1671E4426DD1EEE1F479265EBB930838CC38183988235C58EF083097D572910C70F4EF45DC85D7BDD9BBF179A1991E7B9C6ED5C250C19C0C95E2C8AC592B91178549EBCDC6457337398EE90EBE8EF74AE489C0F292BC7E2E5C069287C009CA074C830558EB7C28B88D5D9DA8173EEF59758276B7754E94E588220211ED6DAF4FACB479F08F072860E8FD3847C3528941DFDD3DF243859B273AD437F46B8E0BDA4995F4A8F4E0213BE6C01D14AF030BD348A497588C2FBDA403DB2C2128D95A694002B8D8BB99BD76E8D9A83ACFA8EA10901C8ED8EABA13E6AB987EB492BEB24F1DE90AD09CB3512046A6616DE5105E421A884D2EF6ABE8781196C9E1B048928AB2B36A8EC3218CB989A5A011F0D5037E91B742FE2D858F938A3A061A72A8D57A15D291142B56AC7100F092028C3A0A9D001A5115C18803FDB3BBED5F9BC50AA8BA6E8AF302DCF5606C319058BA33915F81D2AB16829AC833E6FE8B9ACE289D5E6B9C4256835A212BCC099D058077896790372F17FB249E25C6B15F6AE876FA31A0493D926EEC95430C4B16CF124E013080369D91C5F7E6A1B1AD08B6100837F5E0295E97715DE054B902EFE0A04D034DC8787709833C0B0364DBA5FCFBEA92D2A18AFDFE989AAE00EC9AF6C2D37D23729F55E93BACA9CD3539EA3B4C8B011B322477AC1DA54D0F4042FA674D944373171FB8047F7847DE44E714083E9DC850FA0D7BD8BDBCE5FA4E0BDC356F61146042CCA3809B424C70C6821601D218CC61B3F80943297BA9DC412B26D3B2CB76E5436EE63186DCF78402E8B7CD7E310BDB5E2FCF9AA6472E0E3933E8561AE5A7EBE9EA4DD14F720588F69763B8B3417643F1EE536DE7FA9678ECA1B0BCD7685E5EA26C07D38628FF7CA45CED0EF8004B41E6461E1EA61C2B3F20DA8E33272E8DBBE09A7374427301CF432B77B6'
	},
]
