// Copyright © 2024 blackshirt.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
//
// The main SLH-DSA Signature signing testing module
module pslhdsa

import encoding.hex

// Test 1
// Test basic signing and verification
fn test_sign_verify_internal_basic() ! {
	sk := slh_keygen(new_context(.sha2_128f))!
	pk := sk.pubkey()

	msg := 'hello'.bytes()
	addrnd := []u8{len: 12, init: 0x0f}
	sig := slh_sign_internal(msg, sk, addrnd)!

	verified := slh_verify_internal(msg, sig, pk)!
	assert verified == true
}

// Test 2
struct SignShake128fTest {
	sk        string
	pk        string
	message   string
	context   string
	signature string
}

// The test material was adapted from golang version of slh-dsa
fn test_deterministic_sign_verify_shake128f() ! {
	item := SignShake128fTest{
		sk:        '6c1f4a3889984abd0d30e9454e8ae15d423be3aa1b0024599639b0bfb9c41e9fff34692100a04a8e9bea7ab80e2eaf8031e099f8dbdd09e71adf94836e3350b1'
		pk:        'ff34692100a04a8e9bea7ab80e2eaf8031e099f8dbdd09e71adf94836e3350b1'
		message:   '74657374206d657373616765'
		context:   '7465737420636f6e74657874'
		signature: 'fe9a71dc6a6920b113a168b78fdf75e0c33edb3d7302227abc8ed4c4c71def4b2b1ed071eb57129ab6387b43e2ddd659454eb1039fbc61b00dcdc0babaa844bad98628ccc862de4e969b6457ff21fd4cf538a50b89e4b7d77a1554ba16137a4c566e0e5d450876f2dfc4f90b18a578cffeaaad93064f8a5bed56e6a5d98e477253c133899c42eec2896e025f3fffe92f5148ef7875345c223f4fe8a6bad0a50717553037e103acf0d12d0dfd3fa71d30ca2bbc0253ce4d01fbad2002dac53fa029e2c0cc9e9f551e737646d63921aed8558862005b06793a8ebbcb099cfdd83827a4314ec6587485ecc3d93062e93be2d78039e6ca9bc03b12c1562fee0bd2e5cdc7a5614922b8f9bad9ae65f8889db82ae7f5ecb67c34289eed5c34abc8784b797725c07b219dc54cd9991031cd802b84c2b9e0429feff755c1ab380d79e0c7f7bec55db87d5c18517d75f0b2866da80f6b61b07f7394c56486ba1e1da16798f909441158e2589afb2f72a23321e793266573e1328d11fc26ca792de5402e1f6de8615832344a7779f72555448e3ad3795cf448d09d74ba56de6c364f14a6ea3cbacbbdc2a41751e0d213859f9f74e3a78e98afc4df9a04eee68fe86031c101ed43dc32d9ddb85011c04cddd298134faef2c11e0aece865f497c88335741e8a85e5866c2473eb27f9c9a090e79ab49dada78fca2faf3a85b2572a5866ae4ff224c8451920198c04a5d984caf225efce8bbab7dd7967a2719bf22f89529deeb38fb8f880cfb2fd2d2ce3f7ae433260f7bdb78ad78d4f3f506d07a4febf95a7b5ad431081c88b030e9869107a6eb5526c871eae188bbb6428e067150d504ed508b3bf11f0e61f01b11ec0ab26de6e75cfc2ab92b7fea9d3763b4bea54c984c18daa5a3974d9bb93454a318a9193e9e1cf7d24679449dc2d40b11fbdb58bd46c4e3e572b6bde4380570c58fbb12d4bb7c2fb60a7911e8d336e16c55d56c083f69c64de8ec1bcc4bb1b2d09d8af9de23ff6c39ca53471e93f152bc5e51d59edbd6e5546666519f5153e3efe621717c42c96a20876eccd3f93f7a82fbf6595a7af2a57754762bbd31936db4c77d54362d15f37eb7cd72e7ddd940792b3992bff15f81c28a8b1dafa34e217b5bb407f9f16fe2363cd8f063f8548b35cb123d06615133f1672448bc3131b7c5dd5607975dd3960925fa02e984ab4df6cca56b5e24f1b5939621b7777fc919168948769eb912fa160ec1cfbe8284b4c57a59bd9921bb0666a95d5379f59a70b8d232e5c055d9251a90029b9a8cb75a32f54297ae5b4d0c0e7bfdd2a202d65dd52052efa43f60c795c898ac8e6852caba5a8304cc814af44a8bfc97e59043d2487a9724a7a209feddb490ddf17cdc5ea58fa4759e912adcddfc0c43b8a050fd143a2dfdc7f4f9293630792455a03af832212cf82bec2979c89887da4f5f211e8638b7b6eeaf5ea4a22cc72fcd83629215a325f4930027e6584db476269ad47da2948ea3ca87e856a442cb2a4bef2b59b208965d4c5bedb3d8bd10a608b13ef1eb9c06438a2a16b8fe6ea9e35cc346591e3199de6581b5cf81883f82a010614cf52579823a802d2981ee13689b3b29412133a6b7c18030007da842af81f510754468fe90b0b2a2dff44a186104669432dd793bae29ea1793966c43438d4b190d414ccd0d4455c837c55d694308dfd53403bb0cc4b255f56d9329cab21ad44a72f5e5d02fa939c59b5787f3ccd503e95eaa8141387b6d55ea6fd87b519f8caa146a4e60a7071645f3344a3b1af79c4f28367c9120738b4d91945899d958353be4a84a73849e268399a905202e5e3947fde7aa7fd7266222f579a1140f4b5f412b18a7c6e6404eaca3eca437d2bd9723f405eb4f36947539696e6e0901475c99e26b540a3845101125dc1f6d9673d432a48b70344dda574b155c6fc098d241b657c508b45e6a0ea7d8cc79e80fa03f0d24452c63b4bfa90db6e85dbd38c5fd7c09236a8f20a46045216907a14743e638afe760de17542d6d4b2bd121ac1aeb836d3642f403998beb65f865ab9a6fcaa6d0906be63ff0e6b15f387e5c5ceff8ea4d23e06491bdf7dfe3d24264ae9afdc3e25ac8b3362a2c2c4e0ae9fbdabb209f4b04371912864d486a6a000a88ebea1e01b8a6ce96af157fbb8393672d0b8d9e629f9c6c40145ec66dd118a56805919aff3aa96dacd44a3a2bf9160b28ad15fc69ef89da0116a514f05a72a9b98811f6fc9b08214464e3d053a92fad9b7c3a2b9ba10301a81b561c7028f61e222cd2da7e87abd4196b0ac45706d62400fb2c8f0f9b153ccdbc47ac6f0c74d50e276c3820b40355ce90800692b700c59dfce9a410279bf63c29ddf9e673a36e199804e64ac1f494b8e65a1403da48acae189fd4685a245da10d41786234f3b12a11d7e3dd432ba1ad3f084cf45eeeec8a3b5d8991110a34949eb861118d25e3f06c0032bb233da15004db519042e62c359401c7e832534dd912d8b261ae255a5390d85f40bc4e3ecd4eef091aeb9b15b5f4f0c0e02d2c00db095e3c5d3c57275e45ea41d37fcab6f04d807ca96c90c26d7d0c7c2d691dc1870944d9226ff8efa143bc8d48be6ff438e951d21841df58f91fde297b07cba4b193c6d93aa92a4044e886bcaf4bdaf7b3dddb80f348018c9e55fcda8d86372b0da9d219034b635aaf15d711b62ce4bbe30a8216239f80db0a9ab3bdfd6e2f022c36798d72ef6467731a657d5e511c3234f9dfa6db158506f5599eb82dcb79375caea8ce3e786a901bf791602ecef231dcc07a7ed34d346e8581b5dbea796e70bad5c25135a73d1e89b4264f7333a2859b348261d19cdd0b1c6d7aa5cb65d79dbd6618f1fa11a65621af049a30c855066385c4632f9f51b3b4aed9107f395da9adc3bcd2b0c19a6d0ddb1835616a5cc97a1d31d25b8dcdfb68956d79120129c31c3486258ab7d8e36f15581d1138831a5d6be2dbaeeb9c9dcf7b86fa16a75902658650a6c5e81b400dad0666efbd04c2de45b910e73eef4669a142999cc6aa4bb79666b8ec686a38a85be7bcecf9de5580c78b621f752eb7b0e1dd11348d4f4024f3383121c968fc8fc05d692c2dc586b3c0dc47246143cbcdee6a1fa16552decb60466b40dfedb44133673fabc16d8466a7289db3cd5132b3bd14979d5ae8dc8ac54c6d759d608236721cf0deb8b9f73d68f77f58e39b41c351f32eef7d5804695dae1fd87d27ed1254803884de5049e1fa6ce734b894adb08b3ef5b619b18a298426dd6e17665413bbf8040346028a29c8e975d574396ae898985337716db8b87e52de80fc8102996f83652428917ff6ffb399e84b76c991dc892882e33bf34dfb0ed84912cee27a33995ab069bc9d4468944dde805d30934aa1dcbfe434716ea02faffeda9f0b7df083d0a738bd3a96b45a1c5bed586c19127ebe1abe752ed2aa6252c1afe271fe2313937aab2b98243915a170aad8e00fdfa52af16f6bebb2617bfadd09cdf06d07695a8cd0d76e1dfcccc86a83e9510a16d5a6f724262204c5c199d763d96ef9a134167179adf6e09af580fb2a76753ac0197ae096c53dcbd2b388c64c4cd7f5158d93472676766c59a8dee6ebcf6ca8b3744be790b51c4b199a8012ed76357e4fa5a4d869dcd66ff974af5efe252862c528bdf669ebf059edfd57c4923ac141a9cd1657406be03c73303366260723fa5edd76f57a467693b9d68c8cac60177a7a40b5e21006e3bbde28e0a18454a01758c7f0aa5f476e03e71589168047c5553560747711de041eb9f8720b3fcf302d63be4e6b7a7c863dab7e3cf3d70c3c6c0270bb723a795f53e0ab771713cb441d659825a347882acc9b713eee2b6e6d01ee3d7b0152196f4cf6d1550f1d6770f2766c60dda1ceaf5b2fe21f1da674451eb15b8b58544627d9f057fcc5285d163c1648b7dbc6889cb653836071bd4b2e580dfce825c5e68a58b6468db2324062e1d0ef55e578a8eface3da930fb2cf6bc3e7a5017af6e680a3887981fb851b3e943df4a0584f8e3bfd9be10f16c67c3773654ee8906bbb24c8cba6205b7d87cb234b1f4c253e08129aed111479122d9c3371c43db7a512c8addc516496a85e5583835f4710af40f57d8c6f7908056f99762a34ad838d37ef587cf22ddd821851e193563044c0d38a8f6b2902df7a502dea701e7509c1f59161b662d36cb94feb20700cee15ca5d8b0b5996e20e839e7e3bded536b17ae2b5ea8937a16781daf43dd25d41207151fc42352e5a36d162adaeb69bad5cd954dd02187fb610053dbd04231a6b50a640b7d6fced29709b0b6db45a2e200f5cceb6603d6eeb0068337d5d3dc0f782e12d9e76a074a62b52ae9a3dae80a30ba1cca441322306b7a066a0eb58b4f5662f219d65f3a08ba9ff7301a0b41c986c9ddfb05b3b3ee4154f5bad8def82f1e0794480bf56d6c02582034c8a2d9bc99536ad90fc9dc9f79a8d64c38367793410dbc25d52ff29cae0a51769d686eca8920fd1f9c8d5de9ab426b646c44c5b774dce69837b3bb35a58cadb3a43f1a49d6d5ff3e77f6b01590c42093c624aaae49d93eb601d2636f90d79d2a332e7b8c91f5a9d71017b1278c049403de6e44111da49c19180191dff216780b88c091e011f70682ae73ddc34b92e5379f9d886f01cbcdba858b4c7213289647723165a0719a4e67d12d68686aeae0708ce9afc1eebdd60c46b9e7fef25a8a80d422aa348a88f0ceb82498e04bffad5160d1136c5c8fc8b61cef003dc5e2c80b96b47c81a50315131dbf9990c45186636cc325649f1f4f7ed12d8c78f8e70e1d8afb35a730785a193ee04c67e55b33597632c348acf2d02018105bc2f7bddb3ab9defad388f3d2129fbf4c1d6a4decd361f170661016f3a5266d333541ca2940251e3086a6b6800df89749564b3c5f7b45230cf928da121e7ad347352881690302446ae3642a4de7e728bc3bc5bd52fb1b0f10f39f867e50b8c98554ef7fc03c2c205a8016adc87978255825d1ac67481384c4b06e51c51f8fa98a0c36fdf6b2810086372adf82665d9233b49b7cea6e2439a59c92a9e5b3d1dd9513fd496e73c96990119d0bf6821513b3340057ed491e7b79bdc73292db91d12eefb4e9feab56c6d97e0d01e3dc5c1812d88e1ccea9eba6b460d8e7fffeab1266fdac83921651b3decca35830688746cbd09112f4e326f9dd5175f0de6efd433555b64d0354be64cf192ecbc9d4bf0393b14348ac4d230390bb10c42d617ac650e9c8aed2df1681e919a2a18503de9b629c2271381b2f333b8a216dc189e4ff2a95886d66f1ba7b8f91c8bda8477f1ccb5300c485217197b7bfca06c6cc634904f9c4b706b62d98fd9d48b5850c7488479c1867d3a16869141bfafa5a5b4bcacc2dd1ae49cedb3e34ed9b5b364e3e143674999026c9ea396a78b928897e15f52a4da9f2f5288d1e0d87fe8b5686b9f50741683b47924b6b8a31b9d51c5229fa777700975a314396495cf1af574c49599829f5653a976f004e97f201d3fe0dc08baf1d66f3d77b4620d3c8315e751783b9f493a939d358a5dc4e0a7fb2e516aee0e9f9eb1e89d72492c59c5acfc1687aa943334fb4b545438ca741acae4e6674b37cd2aafe46f4418864e0d2b2e794082dd8b0c8109fcc53a578f098fc734d13794c9faf5696faae36ae2207f9fb7096cdffeb90ead0a309aead73888798f6927ef311b6d97a46ecc95053f7bdac1c087b47a0f96dfb6c87ccf50f30ec3f176ef2bfbb778c63b2bef650d8936561b0bdd9a7bb8d469f30984b0d83a026eaeee2c66cbb9950ffa19abc51f7656fdfc8ceefb5f048ab272b39dcd53148038a38dcfa56dc6664b20b1da9f6cf24c5c1c653b5f89a588d1ac7e3ff0a51001a3433dc2e6fc18dbdb68986db2cf53383ff206293e46d3669b1fe36b11f262ae87595b55b73d6405eb8d4ed47fd716cbfb78ad67bcedb53b78d015c40556ff5ff71b09ca08549a75a0345ccfc113841e6c9dbc717b5674833c3a98e7430e24da32f56d15c0cb0a334f7bcec649aefd38a5187673a9a6f45b7c76208d5acfd40e155ccdd0493592baeaa5f86782e0932a1a3719dbf2622cd44c528d813ba02f65f8baa452b0aedc873d3946ad673dcfc28bcd6ec3e4b20343f8c4218422c49b9ab3c02fb6e6f6a41a761b72a5a5677ce80262379bad22af24eca82de2f647e9c01c4b191838143d02b8eb91d27688a943b84a6e3a6753af07326c20dc1478f2badd45077d215de9ecb412279b1e0f227891c312e81ef4c97fc4487901be11145419a87b54c46a1d8b223fbbc14e2d63496e3128179e63d2b87ebb49c0d4e7b4f6beeb41c918ae4211928f6583a19643d124c381e69f32dfead7c0be82f5ae19f3190a1f8d40dbe60ceca99e9fb9e52528086790c357096a28e555c9e814efe76a8e33025d1c234c52be2193384e4a85f43f9103f4d112947cbe474677cd694fd38b13fa81e5aa7e73057236900d55f0c4dc198f1cfb17c81ebe94c326718503a2f0d92ccabc82baacac51879d246f5da24de41b55a8389f1a97dec8a86d6223cc806dd2e1bcba10b5e825314f3be029badf3e50049e833d67ee2f82ede029a4aba6107225435bcc542b1430834d1436e90ec99d914f361a621cca6835589700b967e62b387d12db2020734559166a4665bf29b495f8553831a3d0993ef9a74de5b02336cb7ef02d50be77af68145b9446df3472f776916dee44858ec4a93f165a030009cb22fec065e927e191b4c11ec4382dcdbf718b5ff4a456a69bbb77c7bc11fe1a496b739e06be873bd7415993a6f56bdc7c4ccdb9bf05a94d86ae72bfdad0477939c8727c97c4372817267cc8d308d5b6b2ee39a6f8b8a5ced8ef64d3736f003556cf505450f291570a0769840ac8265b674b1b8402c5d9729e940c1b5065c25a06303de6a98e0103d75ce6b9113144996572776baea1012c94f77bc02c0ad0b66df9b84e2afe066a79666123945e70f4bfc71c6693bef499f370c596059e6644da70c024faeb837f22cca4cd79732be51f44c524f73318fe5b58b1d5002025bb09d8b0dc6bf3dc74a65eebdb7f4e6eb11c2fc5c7f4e6aae121752d456b58da560dc73fa4e0ba64f4951636202ea53aaa4c638dc25a8c95ab8a21f3236e5f9b651e1287b1b775ca6a80f97723490dfa606937b0194b250e450149aa4f3bb961bd9ddfea2d43ec5983ea8907d5b96b09644e9e33669a6c3f5e2760379ac33949976915ebd25b42a0a9047a8a508079322f40ebf139ef2518c3e8249103792c38406a27bf350ac8f587fd4281961c23266d01d47b583971bc21dff0753fe61f577c38293a8946f7707ac469ac3e6600ae63e7c00e0aa61c5d5013a249e2d3aefc526409b605f86b2ab03bd221770d1196458b8c2683bb9a6189219628349c6aaf184b4131b8e6cdcaec4fb35be9a40ee76b7e184f85278eb69b594140589f360f5d46d87952d0928512a8f39f5cf66705c3347fae879a638a07cbe3da6c71fd51581e2c47ba17ebd2e709243392d1ce6080c91dccc1231d250ccfa44775078fa3886e624418904ec33e434129074065d3b300932425c8133e07b7952b25e92fc4a0e218492c9c7b2af86d4f8cb0f0cf73319a883c253d5899432cd53d8f45422ef202cb863b73247191b07d49c0a2f54354b723bfa2d1aa9ef1e5a7e61e6c0fb82ccf9e34fcf6e1fa9abc55a2dc5f914565b6e20eeb753dc6702bd580aa18013bcc44f6394773858729640b505593acad07f066c194f989362c64bbde6da9ffe6960fabced2d1168d38211969a857f5c26f4c29def3ac031182e7559209dcd14db355fb39a86ab92bcc7f18457ca43c4cffb69f2f6bc269dc09dd40205fa4fb9cbc677e4434b042217cf4fec31d70221e83ffeb0195191ac0c1cb95e908a0cfcc2a6c59be35538b3ead89eb873c4291d241bcd1d1c37bbb1a31a0ffec4be6304ce2dcfd3350905a84fbc4b89bc0aaf2498b4eb27bf92b6efa62bb6404f783a1948d92526a0adb79838a092371278ae6127fd00160cbc3cd90742245d2301520a7253dacbdc814b174cc45dc20b11cbc32448fc4b0778577b966c585fc2d442a0d94fd7c4bc93fe02e39cf52d0f5c2c74b13071af50d380335a0c0df2de60a870bb469b026ed803df0704d79471839b13b0692cb181ba92dd154c56d377aad809b608926a92a92d26db4b2e787c6d71df47123b7d9c37143e6b085ad9fd147a0177814021410b5ef0c13cb481650925c230c273cad81e1049c78297cc0a80d10f1398a5e7dd81e3d84ec3b29e2c6c9871fff71751aa5544c89be541adb5008d0413de11abbc2e290a991969ebe7272daf4664fbf53df9e74f26d925f381caa7d8d9829415aa085b66158f5f7304a0cb035c1b8059c26ab8e6cf78f24bd01a5ed33ff7747055bc8674c1f0ed7863d863b3b6132557b2f165bdd43e9f6cbae8bda6d6cf415491f383b48abeaf1f701639838ba92baa4db96c9340de14fff4bec2fb597f57afbd60347f6bb9f45eef4c0e99f0931de29556a8c8ce75d8d57cc7128917f61506975a9ebee1883b974d0f07533486b2ccd1e13887626a76a7f69a30083956273def434608c1916d5c227a536c527b10c9d0c746753f358c50ef559153fe51da7c394a47581ad17b1eacc06f95e62bf0f370a7cb7446aa6b4498b3d0690426a55a74012517b6843077088898854e042e2775c5eb6da339ab00657e79205a6f0d647b5ea7ab147f1bd680b37e27504e6fa213f7f4a4fc6211fdcc4eebe820d03e7e508a52575ccf1891d999d65f33bbfadc8c089539b0b266b4058f51aad4d982b267c27d5d3346fc2075ddcfa280752b1456e7b036fa5b917b1f17f07ae62c6b17fd22cc5c5d45e1dd204eb5e9c68af73ae6440a1e022eba2d1ee762f5c74dd9a83ed084a3aa4abad10e8f99be21da0e4bcd4aa24cea11ccdd1c245128091de51eb1f9055febf0f8894a0d82952d22efeb35a588a310e8b97e25e08cc41cec02f45d0d807ae45b80c6b3f353f0edbb79a489edbc3713ca011c8e75834570219ea410a89930ac9693bc4df70ae440c0eda82971b25ff34844798f2ffb82841033fbed47f4d8a580180a02c9ef204f4fe4419526af630aff0dea380c672aed4eb512d44af696618c3167b893cdf8663e9e201003e09e08ceba90dd3bbd2947d1e8d0797308112630c24a5396dc90d68dba816cb36dd930d6b527d787cc422819e40cf546cd8cd4ce688f77d19793885967e9c3b62a998fd691c4c5c1a2b6cf670e440fcf0fd36a56ff0f6488a925cb01d6fa661fd76ebadbfcdbab392230bf0a455c479572b74f4361850fd63fd9c7b3229d1b6615ec6c39a6c50af63d008c2786086b9788a675330f415b646de2859a5a11b1d375296221147a7d1d6f47c7aa61b43b61a6007c1a6bafc672bf1bd060f589dc8c6d0cf2891de0ace3a89a32c15587425a1a73ca1ffe6b90a51fb90b6c0a0bfb70e01f2c397ecf9352d8a9b4ae7a51f9aadf6d69c54c642b5918756fb44fe828778891f5ea5b2d6298c17af6d137f2c4230c96bc2650c040a729000ddee8d097346b9609b21fc81f664b11fc7cab7d9e6d56888a9d7415cb008c71d2c9c307ef74c3e88c52f2676170497f215797577b056e21e879ae21f9a466f647af365746d5da9104a7460423e8f549242e225e0cc05755db25968d5c968dc40788c9c0655f50a0c110cac690eb1f3a414244c17894005e2d1ff8f3cfb9e080cce53b4ca6d79113adf81d5120064666d1940b4ded5597a0f829582e407efaf079f7315d18c8577cdf6908bd376907917470c27d053dd533848b18f6497fa1c438b8f486e465f25f23fda2ff57f92157baea16d57d6194fae43d01f26b8caef9d11b4f65138226c3d5f8260edf1648ca82e60af4f83145d9fbb9b815539987f66ea433ac134606fcfbbaa7d2fc16958467a682bf36e1d729880af6f0301625d36971949bc964c54728542609a8180f277f8be971a11ca0c975b3d49c2b8326a9cf1365cfd939fd6fe5942bc9ba42e88c449d67fdfa02722373fd711ab43caec386cf8f64f239cc24de3ed85b896d2c3e35e35a2770ef648cafa00dc4528337f59a3050d76387af977109feaf23921c500a342f07587913f48b0ccd9e592e33f870f119a34b5011cc0739c0d323f2382e4f4687fd4a561059119b7cfd54ccd904a5d85e8cfa0a763c024d889f1ec84807331ed46e470e3cd82766524a43fffc41395199f3e788532a0d6499a2b2fd80bccb25955fef7d05c32fd7f5d4dfd1d03a353cc0c221cbfbc19b161be9523aa4c9b696d4c3090d6c83f103140da09a29f6343f95c7df927fc3ff98e32ca1061c9cf5b2b71421170ef8fed15097ae55cff63d5272a36ff59be0ae635ee5abc2cf1afabde708df20abf4b93aa66ff5583a2f4c2b258bc3832aa1da9b585442a7e7a1863ed9d91ff7783a0d82a0357c0ebcf72bf4429f98ed5a03a03b429a4a307b84822035b55913eeff303259b4098911ed8a79588eba2922950cbeeff9992661548a51f3f121aee303f44ab5da5d72e4722d076befddccc571aa9114a2e6ec0c426b5ee12c3b9ede8dfb879c6ce0ced9c9fa7d75d9d5a5dfb74e8f08eec199d2d63b140e9a1ca61449eef7472cc548ecbfa56f038a559793dcf1f6299b7192b8179d4b39c0f3a6290d5966e25f12195e0babfe27c550fc3abead9d7bdcbe42572179b8d7571b32e5bfacfcd983c24c962262b006b368ab426e8c41316f1703c20f0f3333a59f3b2e7adc515af6c7d0943a8b7e36bfc516e75bd3653a723f8bd6e93506b62efb3bd4191f4d4e557255f9c5900910304cba2e3762005d47e393ce6cca93743291801584ad5c44c234df4bc6304c9c05a5f25e0799fc7ee9510a4012e6b7961508790993b674eafb5ef508641b39dc91981ada69551ab4e99b747eaf33e047554ec8d08890114c6a123787a41228455c3f8d5ddcc81cecaee7814337370c26436862fd1fcb67d61b27c39da5a22c8eaa3946df767d93f5c2a7f271fc10dc389c2891c7aa9ad9b26b029cd4995906a8a2e09948ffee512569f4f7a7567dff3693ba809ad7c6b65b31227ffeb247feb5fa5776b302c9b5a2b0f0b2369e0ced87a95849a10bbd075dec78f031f3bfc61e52e85c64633e2d98fcbcaf46a8a808bd474d2ff844fcab695c4f30dd530bdbafc336e6e71ec454ffa46d450dd138ce9cdaafc3f4492f60083a2b39b92aeb452cede7ee34376ee49522272180c4bbeec208dc3e23363328d0be9f6cb219455784fca3aa79b9c4a11cc84ba08ecef032c9cee34804f8f9031c247e23bd60c362484b90b22682c328d7efbfb6489db36e5fe8f3a8a2e65bb22415606f3f0507c7953509846f5d4cc4ac52d1b320d791541542e1a0611224b5fbb4e5f812047adb6609d2f0a933dfb1a44894f8efcd8a73bb1bf2dcd1f2554b92ff587077023fe5152b8a6d3f542fa55f9ecded7c785e968de0ac10e92ebd5d0ccc76dcc1cbb2d8cf0c7b9891e65d0594cca8074bde24efdca6a1ae6f5e738ddf78c57087ac30540ee745a10bc50439e5654487cd1dda7739640456d0fca1b2cf5371fb8a05f628115de0ac8b3fbbfc6295c7a9d15caf91804766e7cb3ab2598f4027940b1199e17667f6b171698e76231ee4f379210a61c15a195e5bf958f6ce6d06845bf725c854e7f65f1132463676618cd3d671dedb0c454db2f17392f77546206a016a9ba3239ee98c9085b2504df3103454cc1d7d8adc86d687bf9bed0b22163c599b3a97ce5d5397739734aad2a3ea59268c6092647a6b597b41265bd7e8c3812dd0e20b3318da3e0cfc86392d2bbd32f86642407b932a9831184501806a79f3e5ba903f5b9616e515d8a481cf002b2b80ca61ad25ce5f6e31fd2f98f85d40d665b499f0ab5b8447e491ef047a011cc3ca49449b435c7eb170f380342065430934530515a88ca6a7e26a0100d8dd4af6c69176ad2c43cb4094923fee5c0c06f356820925d4277c8aed69e4746292227034896864ab586895ee376004e264b71105df14622daeffb2951f4298d2a99b61d4a5237a2878b7b05060f4071455b2986805822052ce163b6aafd8e944c62f4174f3847d7c4911e1b6343c91a06462e05e02cc32a0a519ba99f8dcb7dcad2630ad7d6a75857629c56adcdc218212589a67712bec8608242acc154f0c9ef76e63b1b975e4c23f49e4f86ae9853be20db68b453eb32931d4ff500f2b099667ddeffffbf4ccd020f51b26725a1d87a735e9794436b446d51be75b5d98c707b1376aebad8d1f12ac3b842e81362afbb075af11f5271e254de0d13dd4bc538af2a5f15047ed62269184abd61129a464faf245917c491fd6f343fb19a6a4e1dc4c87f71d9bf81275568a2376b7c2bd12b2e6a4cc5776add167a2c6156ac02b24d0d7952e41b180a14ed43b49e40aa4de12bd32725027e10c5315983bcc36f7a777db224f57da964b959969b6f34eec76e962a08141a0251b05ba7a14b9a252bb8e9cbc603338bab442e5c9efc9025a79d22482bd3b0f832ebc27648f58636e3d2bad63c1b9f399e90d9c82d4a1be5cf55bbd8ad0718cac5ad70565aa5dd623f9a09038ff7bb748f6e9a4e76aa969b92dcdf5d6d422e254a30562370cb86c36fd2662441681734a5136db2ce486ed7d2e5df55f403b46ccddcf85d023dd9f5642b56dba9bc406078f9a77dbbecd6d1da4d4534da6dbcc50e754e06fae8efb584c1ca302484532c8b6ffcba8365a80b05bcf5e37efe9f7b18a7e3c89e5d4d31d81a75722eded4cf94e57d41c6825f7433b414ab599d93bf1efda78fe5bdf431c6340ec8ff46f1be76a23d25bd3238706ac1db6116483332bec7b5c68597a8543b50754a8be30a2190dd80d4ecaf821bfce9745e3e994f84a5ef28a791597fe0354eacc0b93c0cd003671de34f2b4aa5d709d2552cc4cfdeeb9ba55e8cb451a4aade229ea03809bbe754ca56b51865582c7b16fc55b51eed9143ec1ff44a395010fe19ed4b0634856403908b5f29883c4f84cec33af1c776335f5b2d27df7045a01ee833519d8ecb27dc7c356d6a311f92f06614cb25960ef6a74ab7ccebc2202c88b530a00a6db036c33b44d75ca47e697ac73cba8d8691da6083a0551984ff73c3456a6a54cc54b280d99c3069ae0ce3f02df6b25c4f6298920ae3262c69589c89f19acae4f57d9966a560082021091ba55162eab845bea4d421dc15ab2e4a48272b4a3a402190fa758e49aa9c9ad56c19b94ed8b66cadc26e79a281d1951d943af73837d599c55862091e459c9b8722c96c13b32637dd6729a422d5725dc75866c0a1773e249876b3cc2a867645b8325d67fcb4716e3422c93bf4e56cb2ca692d44866eb2b749e15070d91803747c80c6dfde7705ca6f60087898ca6e84d7771396ca850b01ddd3c7ed2841cb95e295e0dad6bf1ad07f740868c9792191d5364ecccbaa497517ceda3eda2d6e3098f469988bacb6498e0a3a0d180ba63c385f30098766a18d5c208c67e7bb5151cb81c880d6cab5b56bc382c03984a849a6b1080683136e829886e1e4da235fca9c69ea6705f15e253aabae1d5713569ede6219031effb5104e98bc54024e5803f316f6f8f7c7f4b9506ca9614925d532c0fada5c8aa1a6cb98a609aaa8dc75c539790a9688a06deb15d42781ce0e19ef86071a5422bd716ac4621971b9d18fe0b029709d203369a8b2cf91793fd0e5c874e2054516493a2f5aaa9b08feec28a99e9a86f70ee814bf64dc0d02c0c23e7b6117f56ccdefd72e846fa8194c697758eb2e39c0007651b0910e286f98866d006a7f0f1daa037b8370d0600ba4b5dbcc3a3ee25ca3ff65037ae9d823c71483c67dbadc687e6135735913db2e2cb2697efc8429959947b11c227976fe6ea4ef17b4cb6882ce49d5385acf1a7444bbe4048f5d8a97d2fcab42987048541e183bacaadd9d82b01bbbdf2379891ae6ad6414d81df34029ace237aba81cc873c9adbdb3f698899b7875751f111984c679d1be6baa0bc79f0401eaadb1d13da3cebf7da05362502b150d9525c2061381d6bf024b91487b616cfd27734f0bfe58bee3ad578882e70e0036aa1699a49a9cfd1d6768d548cf771236c3925c9840fbf960eedcb19346ebf9aa97c47b9f88e74590026e5fa0a492835f358a8bc0611d9b9130ab8ecd99059a4d5eb35a18e9be0785e316050c3480c9efb480b21c530b01e94fcbdb1704ac0f2a4feb547a32048b9c5a3dd405aebad03d9f13004a853d8cadfaf12fdd84c636b7f237754f5a4899e93fe4b531b9e0cbb6edb4c25fea316ea729cd710f049fc1aff1d3348ec0c30c53835cc49b2a022d9e3153b4d5c0a2bab84e17b40fcc2384b7cee7283c332f5e751b1162c1f8f5aecaa80fb8b0999785ac49c9096fcdb264884e8e00afa799b23bd69fb3800cc5558c33f2aa88218a9197cf5feb9ee3b27a64c5e32b5dde67955e8497e3b429dfef1f4c29990feecf9b00f0f32f818cf789f89d03f49c90a12246bc895531fac453ed92f4d4df1c1a27d829a574b3827d12385b4ed4da1e5e537494e9a929ba58858ab602e6cb36b5d82ea2756c2c204a605cfafeabd61c729a9487a70b05b63d2a55883ad4b7f62f67ab29b85e7a5ed25605614ebccfd423eff83b1386102990feda815c0e5fdc9c44e440948e93d0d42519f0dba3b62430f2c5a7d595a3e09f2e0388dff86515ec45bb10593990e769e7731dcf203a82559ce526fb9478f7afa201ec6b3abe946f4453aa0c3447b1d0d512bc0739b2959b2e7e58c67dcae6a84da2c8ccafc9538a4691f33ceec74f4992ef451a5a66d11315162fa6378d796ccd498f44454fed63c9d7bb7402c76eea5728330ca929ab87a622114b205f8b6ff871e18888ab95edb4c5078393c5f6faf34ddaed97f445c142c96604bcca4e100f9ad7f79e96e3c4ae17f4f7caf8b1c28c152ffe520c36bf8073c4ecfe5057b9af45dc37fcfddc633e9b29eaff7dd2ed16783555d2e07c718eb418b805d631ad2393dc06dc385481b2554c27001f14a13886a3aefb430ca0ff0ae88a8050773c04b57a1498d066f8e067ccba6db31f43ea450cd05b5b5a5ad1202e77c006e6b399b7fd09bc7f5019965f4e7de2f86abf023301aea538046689a3a2e3f7c862fc364f96fe704a70ecf267ee7367bc66ac3b06e9079e269c2586028817c4ddf092e11a2f0400dd3e08a8588f24b1865ee2eddeac65793d6dfef5157f4d934650fc938c6f77ca440d689b6c76f23544f89ba7562439de0991c2bc98d218209ff06d40f7e02bf8af6b60259b6f2da43c0349b518c2847f0954f800a009964549795e0feaa5b219073ffa4045ec1c1973fdba8f4abdaa07af742ed4d9057ddabdfe07d1d6d5820f519b5c33c7271f71699a90459337bafc610e259d2c41b6b88610ec390fe69976e905eb53d6585af86b7a09abe453d87fca735d6701d84d129a1735d57b94104759eefe094773d8c2aa3b6355c8f2abfdd88870eb030b4ccfed7e60caade345c073baeb7d8ff6244cab6aab68b1b23c22569ea109273511d3603549532733b4a29c5f3f3b9d2c74cbe1e24d78a38aa499d6dec331e2853737bc0469221da2caad2a993e66358db514eb0b464ace04db7836534d79da5b083ce323a03f0ac08772ca7150709f5c0f0781b90e0635ee4b3e10a9c97b3e56a697a7ad60b46fd843ef9c47c42838de063b485828a746d23feb5fe9ced53246f5c68954e6d61d7c0565b0326d9f5a31d892031fe838eb0951403862956409e24a5d40c7d5217ef4ecabf4c44ae33e2685e03ae70aa29da511df4ea2e45118b0cfb2e2b7d423a2cbb313c1daa5c7901aabd9db1e1939d2fb61c65e7c923436c8193401afe4d114ed481ce308e4ce342830396fee37dc8c8ea876b3a09afb64936415771c5658a2e965f650079efb4d1831f70ebad7ffdf76972dace238d9c527507c10253c55ade027ab8af3a19060eba34880c44a0131586f6b89fc9a269d08e4ed4debf500d39e2da63784ef58d0c3130c55e1001befc3d1bacf503de5d9d6ea5dc0ecf0a776770c45e3ecd515abb16702b8024512ded6d7852cada0a4ae56311bdfc2469abfe624ad337eb113c8b72054805ff5aeb8fc37afeedf6236a641e8ec65cc6607529e5df2f357502e7515a0693d062fac077eb05e5583f8a042b4d919b58520d7bdfbe8c041c3d61d395ca21c5801765797b5cd277e7e3e6f6a3667bfd54b3188645c4b32fd224f6533c3bb2e849522ee224cad226fc54819040da2e558f78a1336118d83baf025ba0fcfee0b90d198a05edf2bb235d1bbf2ab88a73140b841ea6c8591cf9bdecacfb4c48c267b03a0a58521c8048f5f365fe353a6a71ef8c85cc331d469eac7e93500126137f960f9baa00d3ab3d99be6ca03fa3a6bb5fd1e1a32a43e9982d8a58d39bd0364154125abc1f252b98bf5a5fb0b170d3c3702ed9c7a0f96bf9e39534359f85257f2ff249305603f16fcc24e66dd441e36cc547bb68b05dc31e5ad0cfb78194943d30d0c3866ee448080a750961967485911259eb3fe8c94adfc7a27ee3ba7bd92689c8fe1e8cb01fe7173d99380d83aee9e2b9647c4e5a7ac76aa3d402ae0d1865025017ffd57880cb3d602a3b02fcb0caafc8dc2c60ebeeb73eb1370cfd5bce4e74330c0c2f2b6eef45963ba1cda096581db0da60764fb61febe5d53fc54010b41bcd2604d2ddba53d6ab79c2fce3e79583426590d78bc512a20cf3ba6d0ed852e5626e8f99c0206d429eefe6a5907f768e0f644fe46ff7e3ddfdcec384a629e1ecc310ccefe22239a56db565e3162200c23a7e1181371e9c42996ce2de53c58458599d171fdb50960e3021e495c91ba619ee5330027dbed107dbf1b6ff7b2f7dbbe74a1e5ab56af39da177452ae16bb966f9ea9c075286647ab4bc37b8c201fda72b3bf4d1d2b6b7f57c3dc95fe5b62383bdf835cfcd541ba49f7d7f3413a81860787bb11a8676949d217cc58a7c6f56895ded636e3931dd35b538e494b58678ffd4292a0b14e19c4c9584ee73dfb9fbf1ebbaa8441b3637d11d4caa316686ea36a9ea9d4117aace27f95acb7e176dd4ba9f6d934c479142fb8c16e7a7c29120f920bca136116b783d31c107932cb784d37f09c13bed947ae4dea7706072cf2f40dd782ed099361e85fad0629f4dfb3b7fcae39719f29755db918c4b76f378e0602593152782ef7b6e09d2ea07d3eab79bad9994f6b3c7c9a6382ec80bce1c089c3eae8b66f6e7b634a6dd60255d38df1af82eeb5a61e37b7d61c4abb065019a311aa6e589e8bb70fefa6083a66ee0d30b9b0fc55fa0bcdfd499e5c37bda3aca12511fb747f836c6afd7404b68fe4fc5e7a51feec40a89f35508dd8ec8f10d22b8ff874de5577699cf5e287b00360987fc7c95997288895417e2fe259852d4db215f6962b7e93039cbaeb598873ac0dbbfaf468217213db3b8537aad4874268652837038a74f05f518e8fc4720b12c3169b2e4f0ce398a485ceabd435ce109a3096b79a0a5e534b0b18b4457e3c0f04f829cb2190901b0036512dc7fdd27a8b45d453c40a1a28b26f46abc04aa17fb47b8dbf52a74b8db1c9bdab2cc4472b975ab46632f881e76a208fa7c30a46f626c25b4fccda548254f9538c7037bf837e68cf467d0802f0659956a197d5cfc6035dd159a1062f1f2b606b9d21dbbff8353cca54cad73f9f20719892c6e6f49eac2e7ac2c7c4d3620393dcf4d7db831fc94e5307c4ad5ba03688ed2ae2191aef1dd38e09dfb84a79b73e6c7a39950075c9fefb71e6e18c700552c4345183d0ea0d227c32bf90c6c9fcd5ff5c63b0f497e8e26c03bd26690b99668656d1c08b923bf95b1a9760c2dbb845aa57641ada383c128f807ae1a19656f98afd6da6d5c03b67ef7fadb40902ba79ae8ad40957e41bc9a0c964995c96c9aa7ee9ad09356ea4cf0f327363bd61d9edc1bee40c3d7b797d44a796a5d45cc7a45add759f9dec33e7c7136cc761df1848a7eb264551e0016bcc4aeb96fe37c64d2ea1be3865e75c4032fee1f554bd128ed832d983de7d7d54e58252dec762224092dde57c08232a61d9fa172aef9be5c7a282f72bf481e44da92e7ee18969ff7d7a770299795704feb238decd53e34f72fe1db61424d8d26567f2004cf7970cc075f9f1212449ee0a1f57a19aa0478e2b9446114ffcd0c3c49036214a60927fac1e45dbed7ddaffee046bf7d7566df98cfebec14497e9dbfdae00193b97255ac28ec425e908a5c969325dc21e91527f60d0a95499c95e6115b3b7fb81f88120a51fbdd6b2d6c6ab6218cf43c73487d4866f7260c778b3570b086b401d5ea852d51e5601d014eb14fd7b87e3add6db645f45e123b8a77c2b6e91cd7690fcbd9a77e64c236dc74ff23b2a4eb49d5a1d9a6b92801f191b0fc055882cbf01fce355bf1850f87018aaddbbb5a27e7dc3fe9f52b9951f360f2fba90d1508ce33987c729cb3028991d9e780687d8b06e9e3149626b5e957466a0fddebf21f71871cab2cccb4cb6df068e1328a16fbe119f262d73943f1d0bd6f93d7e1a03ad0fba0ec719e7e30f909ea1518404d6689e9a08e3aef56f0baa5812728094a1971e4ff57b809a9cc25b0052af506fce69e563f1821d16aa20dc2fe53c25973b1341831671ecb1f480b4fcbe6dab5d3686393377d5d8651d02df0c0a61df373a0778147c1f0dad3372dc0b61f9a1882f74f56dd861249ec011d8ae668830ffa9f71280618d43a468433e9dda9ca3c61843771cd5f72fa1c4a84dfc8890ed1d2942f6eb594d88c2a67978f10f050eb905efae38bcaaa5430c796584c664a4a98d6104fe6dbc853a2f67085c3a5bb917a155ac129937df24e197ea8caac5284e45d4c3435f3c3a5904f0fe264bf4f8d9e2827f04a92b8a8ca828b01d59ebf8c4d12f64af564ea53a9bd93c273118c66a6b7ce4bc145b46df232d1daea41f8ae96701adb148618d9b137eb8b6b32af6abbd593dec821af5ffc6a14fab893556d75260af9ba48e65173f32bab22db4e3790032d7fd249083338bace8ab1bd82c53ec211a3df7bf239b9f602b83ff26e1f2ef0859bdcddf9f3432675751546d5c8d06dd110bc8d63e7c478cfc7d63039e443ccc5fe283f6c60ecfac4bcf61c3e1ca8c837d5f33cece6def60c662d015665d4ff9ca9bdabe55280c721c2fe27e6deffd9387662b00c9a51b7916692d221cb81d29204fda7744cac65b05e911445158061182d123f573f897fd7e48bab6b281e1c8f397e072a573d62cb143dceeab4dc2cef3f1acd50218f72d06dbdc3cdd2186fcf9c753f905f5a6a382fa70d1aa5a59b631b1bfaae7f48a40dc624126c50792129b47fc63ea271deb7f48a1c8e975ab81ce9f3cfca585b63d3a8ae7e46e860aad2aed5664d12df8838d5f1e17154be7e7b8c99d351a061795741024bbea3c506a2c806689418a700447799dc1968d48d8624116342043e3872187628f1349939f5c24cf17c1d4c9dc0af002450aa5a5951bd486c4ebfb90c7aba880e2d1e542bacd9802894d5b2ea4e37c9c5008c83b60ebebb39e294baa3ab87a0bacdc1ebfb98a72b26331ccb69f467689e3d9be5df836c55ca1dc02fab0b54483e62f0b54a98d0176ba794e859975741eebd2cef586371608a7e447a5816fb18e58a69476174b985b5e1a46331be7677d94bb1d3c3f0be201db1f68b7891f50dde37c455d2b4a6464df49f33a027d46ccb1841e5d949e6a45a37c185dc88057d32d4d970f01208a8f6b9148e6d8c054177439653780ade95d4b172e3d63eb03797d0b59a1e77873eee28bec93c1b446b0020309133909f8649d46ca443190733a1389aed61ce8e3f3defcc847ad656b15f051c9966eb04ec8294e61863425dd67f934bcd1f4d73707608eed8691c83c1da29a68d282625c571de2b3e7cac472523de0d93f72af877824dd9ac3b2cf043e6a43c7b4bebe26fc96d695b402018047713ec5691f3c2947a5e13fabbce090794e0557fc267a8453e39d4bca4241609d3b87e27afd399e2318f7b21a70ea1fc4b4f652ddd5ea3cb3a621dc9e88ec6fbc30575909b43fbbb75df06c67be8e545e8caad30d1fcc576acb6941cc2ca08d0255f30788e754d7f486b4f5adc1d2e99a56bfad1038b10ba9eed3173a7f5b67ea5111844893bbc056aed3d024f47693fa8082a6fd42b7889580936a6830c1cc141bc103999249422ec786deb4ee02c2dc78171956da786e82bcd59b83a2039c38c2e5802ff823e31bcd32e0375f3cd7526de586c52698d37e60399d357a4920dae9194fec4c66e19c259df5a2d3e0dd1a103917fea0a2c71560cdae449fc90e12632de6d1c642d4f2d8dc85b32a78d9bd36eec20fd67c0030053ef1dc7ef85713e3c181fc463e97ddd27019fcc387cb7a1097e1111ff7564f20738a0fa25b489bf430efe02c7da1035a78913109c4071bc2644b641fc0643f305154de1f86a13347346d2f7742ddcf2bcf7cd36a3780a1730a03cd0da21aa20a3987c0bb784a9db2dfd7374b4482e1d29111b3121e0cee68c99748c6bb62c32aadce5b540ae453e3e098df888184c192865fc34110ff1eec590e80d8b841e5a124de23c44926978b83a69ff3435927b16c101aeb095251e7ffdefd2b2e417d666b33be6e40e3a25f4b9b932397a486e0220a0bbe65b868e28e0df0ce2b9ad6917e336f0c56b12b822c74bf2e64076bdb19ff49e5090394c9234621512a8348866b0a1dd274d0afb465bb8fac8d7d4951190caa5f7b2efe6f3a2f30df89b9a33f2140dde476d2448191da1d135e2b491699630e72a9fc2166f718ac9a6e607e27fe98e836533d168f2e47695fd08883bba9c536abd38cb0409a55950e1962069b0a0ffedf735dc0ebd7d20b2019a9bb99d325643856b0fa3c5472a3710b202e6a6ca04e1277c4cdb2f08fb28bf3db7f1fae32c4664c6a559a346246c18dd9595b2e2c4467281ec962e6665bf97db482bc28b9eb07868e32ec57fa6e9071b85339cfa1891cd1c3c6d0f8d49803cf3de08aa326e66106fae629b628d54bcecb706b59284aaa565e26070865f2495182903622de0820636720b50c61261f0e3daf28cf6628f3a814cd63eb11ee5a3febcbb6d67f571149e9229dd0958b648f091aac40ec65aaae1b323102d94e186479d86de0e6bd990500e400ead65bc30b263d4e20e51f43779ebc51d421d4482e124d6b53e90bff2e70189b10c9c333357b456c114c014c639b080a79ae0df87745e52a794d38f1549e9f923f910a69bb4d6ed0f621150010c78be831d2c0b2fbe130c6220e9333889ef3b39805d13464b0ba3ea9e480e7450ea0e56686ff8c1a9eb405425d2fc635a8143b8cfa123b73c694c4c1d93d662ef6bd362651cbd650e16225e2f4bc44c258ea9053fc5eaaf5acb542c3f83c4d8e47477e3efdd6562d403bf5345a3b55dd17423307c18ef69ab4bc846e9cca7a51254765fdaf94ae42febd3875a69f2a5ba217e88781c0397089c3367bf1b02223af5284b27f8f57b132a944453e1dbcfce007a68623bbb4e43b79b9a73010dc6fa12678c0058ea1908849ea222941426726732419f3ab91b3c5b408fe7f43629ca360927a7df1bf49c1c1eccc1f30bcc839a86d7e54edca375be862ae1057da12571807e28a118231beb87cfdc8924157f002965208af901a81ce224d7f7bf907b202c5d25b046a4138a72d73a113bfd5af4fbaf226cece8b0a2e9fb7c92764dfeafd41952f283709c2e8a137ba162bdfac3ce88c95b55a2e9c91b84b33df2e437e8082beceeafa3e0745c9e8f714706fd70cb703a945839058e865e99bcc4e666034fafe4d2a86221900eb117f55e40e8e64231330edb62693c63fb95d81a4e6c038b0ccebbfc17d657a168cdd1e9217f460b99a96ce4c2149248decf33201aae98f5b84eaa74f0a8b89dd8953a9a79c12597fcce897ecba29ac79325ec2d12c0534da7a6aeab549265edc354c0837c580c3903f9f99dffa0258c6609fd22a6e69cc044b5f64b0d25a6ade4074393c4875b93a2a16b8638755615c7ba47b6b15a7a3c6b6b499a4d1106e14f079d1423f0dec1e88f9d1f3969b0fc7dcd704c405e071b5064900311cf6b7ba503f46d5df9ccfcd1ffbb5387388dd236f4f9b0379aca1baa4ccca1de8bc232865137e69d28862f91a605c91c911981b4a7141a115b79919a0bc08db928a4ca63f9c4d7225b399a05805d099c4c8a1aa2a069529b9db04834910f9afe9b26b67732472685efe686e63eb8f674a7b8706217c50b9bc27c6c83bfbf5d938c167bab7247f7e692843f3f0c07e098917f9468509f3d8e277c59860a58b1aef288bd9cf2a85c088f9424c0e39d6acf01a0f1e22d91b053526543fc45411f267b93343d26a79616a569cf932215468704315ad1fa8a552afd5907a2e1e6ca80b4f7c589d4f466016d1e8f798f68b92d6a1777173b49c4eaa4a44a48984648c1ffa692411b7f86e0b170aa6720a20d840391d9eaa2e1a9e98712469b4f782e2e1897371892a54f24e2a4b2b4ddd38eafa1ebbf3012f77f08d958d300e038b9a266c43eb85c7bfa06ab7e3ecb509d8ee64d1893bea13ed5a4412d8b9a5f8ffe49f9dacdcae2ec62f0bfccb5f2cf53a79ad586b0606a5c76d3fb7ee7841abb198cc22d939db930d40f66201d42baabb0909f0c812c7bed933bb9ac0d9c3634f3350bde8199ae549a67acbabc49374ef3736fc8dd8bbbe46b4e794e34a1a5d24d150f44a49e6a1f90534a0c9f08343395128d63f7bb57e286a7beb691dc4bfb545301e9d9a50bf864337dd7b225cdee8062420c3b4c7bf80d2faefd46097059b7bdfcb3c9658d71ac4e42ec4a031261f9cfe368d9defd56754b04f5418145de65c1ea84467eeff5f2d7f1132a6aee5e0788d4d1db723f6aa6b428e015b05a5ba9ad2c80e894a0b4fc80f509337905901f33082806122109554fc7700ac34128468d9d9860325eac1219ed811ab7440be24fecc678a91b8475a70756c13df1e7ff04ff260e2b9881ca633d2291e39e204114eea3ab02a845737f3c0dcc71573a0bdcf5a9e3571f7466ad7a1013e18c01e38fdde8084c2282d8131c8e27ac5d5d281f876cc08a5e90fe487d41181a2319d74947271e986b793d578f311d79fe88fe0c60331022261e53b679b3806946a7632e0007ba2fc96066b5d9177f4921c78326edeee1a9132fee1817ba97dd298b8759fa7b6834d4ff463087efdcc29c53e304a12dfd5a57d98c49c2ccb0431794143b2b7f0c718ebd4d98760d3550655a38237d52ab138655cec5c4ba187359cd7c29d83b0011e45dcb659a99dea8be0e9e9d35e8b9eef0cad8eefe3400e10e716676e31b6d30992ecc6f85f774fba7a2a24a2bae0320f1117a2815ea1715bb34604a2c503be13dd215de35c47d4c4d41c1fc5b661e6f3a60b33bf8158b697aa0a8f11cf3c0f9c1e3f789a404fcdf59d4b8edf1f0d96013de8a51149c3f3c2bbd1d4da6397ec7abcd02dd878cbee907016d6b99cab7f2eb2682366ebe8def0c9b9ffd28682ac8b3f25b3dff231e6c5e96a2ffd0112dc5b6a5fde1d2423ac8e309514f71343212586344b143557b6cb9f28dc150ce880c6db8ed830f21a5ca7b77e4c79669bed64bbc7b1240fe2f1d2754235430b9c57f7d7873b1a6128ac4ba8f4286ad7bade497959e57b094c0306b9f3af1077bffa974a82b4ccec032dbe4640ac4dd526b4b66c4415dffd975cf79c0792a124664eb6575539676c5eaba5b918ddb65605de7c5f01a4bf620c7622436c3299d3d5afe66ab92e67847ce07457dd6e130a10463c457ffd67e8563dd27d8ab3b97380a1b2fdbe1f33ffe24307ffba9989ddc2fe053bf477694af974c9b606d4b6e5b2798020c160edbf4976d26ac020670885e575f99b28b3ccb61b04a387f92e219b39d679115bfa1acb700e77151cbff9c6d9c2883439fcab36bc13776472729ba231195822b8a87864286977e3bc076259b837653af945d03f76ccda6dbffe92c4595db461e6bfa6fecb18bce2bcf1c6b543af30c6e4d9c76d5023949ad273158ecc22c7619ef83f21a6b95b9ffc68d0ea60471c6461fb10399ce9d311f13e5df8bdabe0f'
	}

	// Its Shake128f Context
	c := new_context(.shake_128f)

	skb := hex.decode(item.sk)!
	assert skb.len == 4 * c.prm.n

	pkb := hex.decode(item.pk)!
	assert pkb.len == 2 * c.prm.n
	pk := new_pubkey(c, pkb)!

	msg := hex.decode(item.message)!
	cx := hex.decode(item.context)!
	signature := hex.decode(item.signature)!

	seckey := slh_keygen_from_bytes(c, skb)!
	secpk := seckey.pubkey()

	assert seckey.pkseed == pk.seed
	assert secpk.equal(pk)
	assert secpk.bytes() == pkb
	assert seckey.bytes() == skb

	// sign in deterministic way, use pk.seed for optional randomness
	opt_rand := pk.seed.clone()
	msgout := encode_msg_purehash(cx, msg)
	sig := slh_sign_internal(msgout, seckey, opt_rand)!

	assert sig.bytes() == signature // PASS

	// verified := slh_verify(msg []u8, sig &SLHSignature, cx []u8, pk &PubKey) !bool
	verified := slh_verify_sig(msg, sig, cx, pk)!
	assert verified == true

	// the facing public api slh_verify(msg []u8, sig []u8, cx []u8, pk &PubKey) !bool
	verified2 := slh_verify(msg, sig.bytes(), cx, pk)!
	assert verified2 == true

	// Test with SigningKey.sign API
	// sig is deterministic signature
	mut opt := Options{
		deterministic: true
		testing:       true
		// Its pure SLH-DSA hash generation
		msg_encoding: .pure
	}
	sig2 := seckey.sign(msg, cx, opt)!
	assert sig2 == signature
	verified3 := slh_verify(msg, signature, cx, pk)!
	assert verified3 == true

	verified4 := pk.verify(msg, signature, cx, opt)!
	assert verified4 == true
}

// Test for pure and prehash signature generation (and verification)
fn test_pure_prehash_signature_generation_verify() ! {
	for tg in siggen_cases {
		ctx := new_context_from_name(tg.parameterset)!
		// get message encoding mode
		mode := if tg.prehash == 'pure' {
			MsgEncoding.pure
		} else {
			if tg.prehash == 'prehash' { MsgEncoding.pre } else { MsgEncoding.noencode }
		}
		mut opt := Options{
			deterministic: tg.deterministic
			testing:       true
			msg_encoding:  mode
		}
		for t in tg.tests {
			skb := hex.decode(t.sk)!
			pkb := hex.decode(t.pk)!
			msg := hex.decode(t.message)!
			cx := hex.decode(t.context)!
			addrnd := hex.decode(t.additionalrandomness)!
			sig := hex.decode(t.signature)!

			//
			sk := slh_keygen_from_bytes(ctx, skb)!
			pk := new_pubkey(ctx, pkb)!
			assert sk.pubkey().bytes() == pkb
			assert pk.bytes() == pkb
			assert pk.seed == sk.pkseed

			// get hash function when its pre-hashed mode
			if opt.msg_encoding == .pre {
				hfn, _ := name_to_hfunc(t.hashalg)!
				opt.hfunc = hfn
			}

			// Get the randomness value
			opt_rnd := if opt.deterministic {
				pk.seed
			} else {
				addrnd
			}
			opt.entropy = opt_rnd

			// dump(opt)
			// SK.sign(msg []u8, cx []u8, opt Options) API
			signature := sk.sign(msg, cx, opt)!
			assert signature == sig

			// verification path
			// verify(msg []u8, sig []u8, cx []u8, opt Options)
			valid := pk.verify(msg, signature, cx, opt)!
			assert valid
		}
	}
}

struct SiggenGroupItem {
	tgid               int
	testtype           string
	parameterset       string
	deterministic      bool
	signatureinterface string
	prehash            string
	tests              []SiggenCaseItem
}

struct SiggenCaseItem {
	tcid                 int
	deferred             bool
	sk                   string
	pk                   string
	message              string
	context              string
	additionalrandomness string
	hashalg              string
	signature            string
}

const siggen_cases = [
	SiggenGroupItem{
		tgid:               4
		testtype:           'AFT'
		parameterset:       'SLH-DSA-SHA2-192f'
		deterministic:      true
		signatureinterface: 'external'
		prehash:            'prehash'
		tests:              [
			SiggenCaseItem{
				tcid:      27
				deferred:  false
				sk:        '37DEF0C7A10FEF6D26A8131A23489244B9CBB734FBE00FCC802AF9692FC9EE98141A567E56B62C64A4E24346120BE1D916A7525CEEBFA4AF0173B8AB5222A831DC6E5CFB97A39D40A8CC47481A9224A28ABC0D043C65ECEC9C3217FD179B6007'
				pk:        '16A7525CEEBFA4AF0173B8AB5222A831DC6E5CFB97A39D40A8CC47481A9224A28ABC0D043C65ECEC9C3217FD179B6007'
				message:   '96'
				context:   '6E474C49561C210779A79ED515707122BCB941D086EFC6465C186CD079C593A1417689569F3C332AABE3090BA1D904AB16A7253F8C1782F89EEC868946CCEB83B340AF191C87C9E2F9CEE709E76432E2A2B39C644947E1F190A6DE691E2CF892EDF170D3BCA65EB30C6E866D08129E7C55A4B63E5ED87524136CC07B3BD650803CEF1B86E1888658F2FB3DBE6BF55D5021193F6EAC34820878525C42FE50AE492CF2636663BF9695136273E1E1ED766FAFBFCCE91F7D729F567F46771D99BB65DC1EACE1650C0FED035FEC1FD3D887BEC979DCBAB68B67D8D4C97372AC99F4FF8246B969AC40E98B79827587564668CAF1F31111993DAC'
				hashalg:   'SHA2-512/256'
				signature: 'EA7ACC3B71C7E6C9F31BB91645135D63BE0FCA3B2B43865B424568A1445494F2C673E20BE9D367C3939786522EAB7DD5C83C7CB668F7781597B02BD8BB56006278B60E6885CF8B017A24B266126318314CEA3EC7AE1D393A3EFF1410C74781A11FCE2A52CAC52B39AA8A0E5B09537462F68D5B8C056EE7A1105E51E4440C22512882E45A76D3C877DF76935D7158746539D1A5EDD9DB729CAE267C83E729A24DC2368562F515C060B4D1B0332FE563F8A42B96CDD51D2A5042A00E23A49D9CC5E70B0411493C6820D5F64D616249AAD732572849BE8887B98822DFACC71C7D8C7476A857703798676DBB37F9EDEB1509B7F6AE4FF45099660AEE4DA1EFAD791DE267B24D946C44756CF70E7A1FDA3743A37A075BB8994FA1C95AE8D575D8D70AE5AB687A3C3A2F5448D14919943A8D188C81D1C4DE4CDD7FC57A6FFAD6E71D8BC8213FA23C8FF8B4E61BE7E0A96ADA23D53B7F2BBBF8F975A3469594D10C541DDBC72A2071B7DC0EEABDB01A3BF16A7649577D12552450E1EF39894E913F32EED17FC4D3B438E91A5FEA0E91C81C6C1956E8B267321D7D19F17406E0B1647E885B548BCD21A69107BBEDAF7DCE4587D667739E9F1151026E9DB451250AA5313B0CBA0D00F1CBB9AB798B5AB38F9CB7988CA92816D8B2FDEA3F0DBDCD18392C86D12C95022A2157D096B96F0CAC935117CE5A4B991E7CBDF30DB21F1E22FDEC5B99164C4FC9344901E600308B54D7726643BF95932BDC24D3364C8F358755EDE25F23168960C91BC720488D8630A278D5A77D1921CDF9A0C21EF361F188A3A7EB086407C089B4E50ED065E6DFFE300DA0A7BF57FD4469D2B3D2D9FEE893FD86471B2634B14446A158F7E37288E469817DDC3B1327601066AA5AF91056501096768294A1A9E34658D3AA36C4C5F1C0B66DD2B9403C136E9E3ACEE0C4178CF0374D30B081F4629A2F494B240507733C7877E98FD7AC2C32501078E2F6F9F2E48E49FC41F4A63D0EE9B48A5F2A15403B21DF036869C2855F5509B6904EF45C090799E64F4B4C7327D6A7F2AFCE37C85A79FAF06D419F58AFB03ABD08A72838F557D8C9350E7BA541CE4B68FC03344E607D65BAF1E6C3A208715AD9A57DF1A7F9227A56E0DD13AA983E48DB71EEF4D3B82095ED0C5B3F8018094BC839AD282A10CEC80E2FB840D9EA6B6196F2AE3BA2A7F7C8911890522B63FB992A025DFF4A7CD40BC74DB3C412CE5CA0C70D3E0CD19D945CED42C64D17AF5ADFAE74FC1F92B90448AB09117E67440A01E51A026022AF876CAC527027ABF0C8B2023A8303972661DDB17584E523B29C4B9157C42A4A8ADB7A9EA4DE021AF536D51817F24E079398A8068A4000DB2A3AACAD313D10CEE84EEFBB4B9AEBDB4CBCFC1C0203B6597A245F97C23CF19512D43874969120987C657AFEF7E4AAD62C03FEB1DFF39BB564637585B2953C6D08041BA570F78700C02ECAAC94F35BDD3B58BD946086AD61EC53C4FD919627026758EEF831D9C2BDB97EEF3148CBA8981958F87CE26D8AA688C736632AAEDF648D2E8C930042C0CF4BFA63A856AC5A7884E16FEE0AA8CA97AB79C604D913DCDB7EF11CC2C7F9A367FAB991F2477E60ECB1FE226444A44547A1BE9595A695C00D8EFC5A476DB17FEA1D0AEE369DB0B565721288177BEF3EBD6032A789011818B4331A6D56FB548BDA2CE70B5A64F1FCF40C24C1D0E1D58811139ED800CE52ED9BB8EC6CDCF3D90787C27CD29E54C115393AFA76D3174798A375779153CE8E53F6F5EEDB36C4617636DED407096892BB470E93F438C7BECE374A1AAF2E7D41EC89FE7F333F560CAADF7583C698799B672EDD42110FEAFFD7BB2A83EAEA434C1F0E0C186E3021602749B38EDB2FBC8324C1FDDFD2BA2CEB4C6C06ED2F2ED8BDBE423BA62CCE1691C42FE71350DB9B17EA56240436B4BCF9C774E820D4C5C56CBB34AB2FF10A52F06EFE8A30CCA532396AF8B8CFFBA8847F46BA022E84E68369684CC81377082146DDE0117BDF73B4AD213FC907FE649635E9172C3DE3D5DECD286AB66F35D74CE0B86AA020589F4EA49C097547628152BDFD203AC3CFFE3D9AA7825A44384E40A79063FEBAE60884CB0D79BBFDF42F2FA7D9D8D496A9339D4F408A1E636279E8BF80FA3CE2548A3AE609F94E1ED772CDDAE9D46B9514D1BC247BF162037475422A25F3CEDDB2A40E2A77C29E6C8D588FF9D2747F7BADFA2D08A3D00278E753428ACB87695CB5887EEEDC0F34397D5D5A28BF095C3F1773884826F1A9DBA18B99E1AE9B7BC03FC2729F7AD0A5F1E17F95526A333E1AA61E632715B877FA38D2BFF0B5592A97EBE0BBE5B126CEF098FA9C51FC0076677FE284BB899257D1F7A2AD7762A1E3DC0E4D2A55ED09228870DC21101D2445DC0BC5BBDBCC3920BFDA04E8B168ECD36C0AC1441EA9740CB49C3E3D46C5D0F4E783A81C6190957C2E3D805DEAFDD867E04BB0BA56E16B53409271477A8E42C76222DB9E214E7CE03F90F7FB586F1BBB4A8C7ECC2DFAF8B60F0EB044D877A1DCF11D955575AFDEADA0F9A44677FCF774FC255FCECA41AA9088D630E4AC804D36B0FC4D719B3545A243B2950D6AA3DA6ECC223CEDA4170B92B203AF122C17BE5455B4027A97C292C65C587C883BA855C658CE56DB524C190C407587388E6564F5F64E90EF6B4E117B8B7AA13969764F26644029E01A983F472A26B9C3AC1B4E6027767BB7473F41FB9D53C4CEF19AA031688FA42663D77B7493B8DA3176F20225AC80CD5F4DC1828CE8D610FE3F2CF2F53E24662810B54DF1EF5AD43F7C9EF8B83759F7A80076A3B0171C868984C58C0317735CB75DE05CD931A7AD657D126EF1FD601C31D2B2C8C6BF821077174B1C0A6304A4D4D31526845E50CF2C73FDE2727EF7A1CB82264170B54AEF201917CC93896C58AEC59A066111D6927F06E27D64E73C8B439CCC5156EF8061495FD0425175C53CF8AEDD74CECAEB60FB7A6E2BB9649BBCF59BACA235BEF61A48A47D5C66F999EA7050FD148624FB1962E094DCE15F7F863E3C63DDF31F0AF57445EFEBB740C513C3710D0C02C8BF89F359BB53436A053E08C6E2BF4E2AF932D423BA561F83B88E3747556E356B11D9388A7F4E0139973968137E2BE9D9DAAAE55E0D3C7ED0EEEB038C011154DF3F388D002A8BD38382D54C99E8E28E94797C77E3BB16B71C543306D7F4D07A2BBDC6DD7B42A4E7225BF71A87BAB6CC7DD4560ED4C4860B7A9A8D9FABB22AD51A4AFEEC55358C3845B3708FD0EFA1856657FF334A40FB9EE780784469465BE0AC23E4F03C5CA5C53217B3BB89A72BD77452924D84FC05A86461C1549807489B465F0548C759F44AFE14A834FFB3FB267599497395BFB9E5EF29905785FAC95628B75B3FD42AE5B996034CE4298BEC0F41C3E6143E8227BDC79E7CE9CD62849E064EEDDE499251B717472E4C1C6592819FE14BAAA167FADC3B8F868E4ECA00A1C0DA52F479BD24BB621A2795493065B98C2B3B0363EAE743E9763892BD89A352F37320D61618D8120AAA4F32A1C2417E62F3568A0FEC365C0BDF62872797E97145B99F549F5000165B232F855F41DF51F62296AC823E8478AF75A868E47BF878EE612793D386F22E67CCB3C1E4D45A7B4FC7A85AF84D04C61781EF7F7DA6A4845748ABE9E67D2925DE43D17114A80F476F99E06A34B4A213CB8F81537AEC0919608364C3B83740454BEBF85B0763C77C440C34488D3E2CCE1B80AEECE3A3F9EA2C5719154B148E4DFF12AC467AC55B16A0EE4766820BE6ED5510CF38F6C53410C18199151BDDCCCB17B774053CAFBE931856E70E6F4243013AA7283E735790E8BA4D7C809DDD8DFF29C14C8E50745767380D50A9B7A1FF0113C16BCB721CCB0BE3CE981B1BD370651F67AD7AC4838AB432583008DD2B100ADC21E9197841B217D562C7C5859337E279E7F420494036A1608741986B233650A4F2F545702101A24E42665EF347C294FAAFBEC2B7B48C4A6F965DA0AAED9F5D1793C64B1A740480FA02BE4937927CC3839EFA3234F4DC96C1672B650EDB3F6F7ADA3B715E9EAB80BA18D202B71F74827220331372A70C5FA338A5250BCF4511923F991F8C67899512629628B84A7481A3AA5CDD902A416C5739AE707081E9EA38B163DECA6C77F5956A615CD7ADB418F4648831FD3380DD52DA815AC0855FC9D8C5F444C308A1E6CE4617CD8A3036F20F440F53CDC8DD37C4A2ECA03025AD0B9DAEFB6183EB05BC2800D62E10DE579EB9A2C981EEF35EA94D6C8EB3794C7D93AB292E94870FBCB4898624D49358A887A219D4EF51D1CEA3742CFDF5E6C25D11694042A9A7C6038C02F4A79B458BC0DA24ABD41F97EBF31977BC36FAF9450DC610CA59C26CFED862AF87BC39B3A0E5BDDB814D3A82C6FCD5C85908BBFD16F918866D0E52BD9EA957A0D1C9E37998F801DF0F0807BC9CEA5F71BA954FEF1A78EB57142A85F19445C465E71A85DF6D4A20BF0C0AF3EBEFF530DAEA09F3D05C4D4EF1371CD261CAA940FDEC04C7EBAE04613E9561199076CB3049DCB6DA757F4CFFD54BB6FC1F055620826AEF169C9753E23663DD6B142B75C6D48D95329B101CA64309856B8B650B0885D4EFCC9543625A462D66659898D2282E0A7901D8CE98F7EB98FA157050A5C1E2482961997AD805E855DDF3B2815F61953DD88517A9FED37A2FBC9E43A48B26C5D8AC4EA0176FDEA693724EDFDD5D8A4B31782DD0888D246E7CB45D0AA6F40BBE4B0B4A09FE7B156D44847EECB54FDF298C42E41F13D63099BBAAE583EDA33C3944870EF2169D4DD92B9E30D4D69220CA8324BE22FD04A422979726DAC230B23AFE4B0FD127B3572FB620FA1AE38299A681C778F4CFE45A786BA28EC69663F3CD4A3F7B425BC0918C323937D675AC22AFF3FAD3F1ADBD76696E54F7551AC9B5ECEEB1DD9919BF55DFD0951D558A521B692426D7A011C898648420657D3782334D825910609253B2250B056A7F277853AD5D45432F2FE4E05D016E05C7D77F723DF6304EAE4011A12254FD3E22FF9EFE2CD05B947CE8C7FA354D8C39AD289F427A5AB9C389F86A33E75EC59E222EA9B58BA07F4875CDF0A8508E1C4AA03BA266F7740E2B937CF43E6C2D2FD862B993EFE53AAAD53B22621E6B888A9EBD5275CDB1176C2E3C0D2FE0A6D2D942E3F01BDD45B7CF1AC0E43EAFF4C757BA03E82E5DF9697753CD49092380B619E187E1419310F831755CC84A8DAB9EA12547C6DF4E753C36EB3E367C934BB3C76A605EBFB22FAB74F8A290D42F07A23BCB1BBDBA964AEB1576527DDC86ECFAD515881D74C88A9BE03259938E94B95E1814354161166F9B586DC9B144731BC8D758340CA0C3A7A5F09DE0575FE49DE05A6404FBF4490BBAAD1E3F172051E3981825CBB86119B2DF4C8CC8600FD15B913FF90F77C59962815FBC477E4EAD0B0773E12F6B7BE9DC9F011A42BB6F1B70BA226FB2217E6159D0F8CA05FA8BE707206F862E5A9851B88C96DA191823891E75EDC12C4FA3E116F39054388A69609748EEC865E312E2BD63151816EE8DCC3EE32506D1FF504AC385F9EAE2424DFC5E91BE1892158F6C1E5D9CD516BBCC6E542388E82270611E84884C56AEA4881A71D3E26D18687690E1D997C7ED22F6C87A2D9967B973C6932C0C2ADC6F391490F593D3C37FE6E4B5BED92AA5AB0D004049595F4C0EE0E12591CA469E78E3BFED5A3F0706DBA09F6F12E56648A5D9AEB0F55E5C301E6CCA5365AE525E1B419ECF45F17487A46F68A9FA209432F3C08EAF04812D971CEE46012541334130E04AD134EDAD5254FA961EE4186BFA13BFF89E5435600A27F1B4EE7C14BE8E2D999AC9E18B6E02141C865BE1E5B0B14904777E9BE3D46B995151EC34DDCC21934DF62883B6D5EA879CD5C2A1F8246708476F093D591A1D26FBEF53E68D218B63840F44E330ECCC6C3DD08FE0C7B094C0FE784A117C30F651D5C080A40C1E445AA94187AB88A9D91B4CB4A0ED9286D9C1DB994E486A4CC9D51E8F1CC55D6284191B33B84C6C0A800FF279BDA8F9697C55BA78B9D093849BBFA9DBA85B7EAA91956F043443EC1C44CF748A4E48C339E77E58568D4709393B00AEB285B174D6AAB2BD35AC7F2B95064785F6B7C18CD9B0BC13E9BA8A07EAE741DF763C3D3AA8B09B6C3DE1E3A89D0181534812EBE9D364AD783F5C85AAAAD6FAD36EEF025E410073D1FB1E787617CCA17A083BAF14580C0D66ADE71E635BA037CFCBEBAE997565EE60E765805E72D39FAC7C0791B4C258E557F4294B9D9CC882F2AB9377B690A7866172749E9B7D7087C61071273EC0392272A86265FB49408CB6EBC32D260A9A25F73BA3745B8E0C41ECBDC143F61E7FE7955AB86AFAC23507F9E4C935B0F11C55CF6C975AB4F9521FBC82A8AFC2C98C5E7386E6268590E0BA06FAE141274BB9AB5823A7B863E8711743B2D6F3889E782495A99268DDB6BEF2CFB2784D2308834F008014EA5711487E465F3332BF687763A1FEC01DCCEEFC2FD773E433857046A3EE6F9462C0E673F9BC4D9E1E745EF3BA2A9232E01C325BB37BADC7AB9356E338FE1CBA9733AC2F4125346580003E4787329AAAC738DD5695167C0348471793D39D33095D35BAD2AE1532D505479BF8C623B4A629D9230CF750099684C54F9355B3233F3F7DACE92F82123ABA6CAFC3B73E0422F760A5D3B3CD33F4F6277AAA6AC063F756691B9159A65554AD328BE2A5CA1DFF6856069F7C08ABFC381044330DD05D5D7FFE989111E734EF1E64DC04A791E1EDECC0359231850EC3E06E64894871295264D5BB2C784976B7C8C553A3E0D58D6EB4265CF121AB1A543428BC5C87616BD70B491E7B3A18EA4513A5DF033629CB3D26B7A14F00C436A75C372D1B367BFADAFAEF79891B210BDB2159701A9302CCCB309C602CCAE3D8D852025AC3CFBE7738190FC7EC7D439446054A552EB2542317B38BDB993E14372FB3F5B1B61BE40DFEEAA166A4AC2CC6667389A08C3A3469EA673D6A1BAE68BC5688BB3406DAF82166AEB6926D6334DE82F0778B3B632310B3FDAD4E3F039E03CF6C35573E2151DDB9F1F43330B63C82AA8928725B9488CAFD2509173D73D9EBB421D134D5CB851BAD1CF9B397D36E94BD832A239A55EC8E777CDBA67A4AA4E28063D77389033C1981B87EFAD9E2EF11C9EEBB04549EE7537A880E4D53079E88A2E605551B0AC2D221259714C1CA3694595CA675D0A282282CB4DDB73FB0827FDA36319066375EABB6FFE445F52FFD3F2B37D022D3B6B7F650406BD141DC771C682A110202CECC0475ADD0867DA8CCF6D927A537ABC24365B0D2410EFAB0593F3725FBAAB0C7FF2092665FA74257CA8225E4D2CF13F370EDE5CC4FC38C3F0FB06F3DA156AC6FDA17F76CF520106EE4AA7B5CDA30B5DCE0C81C4D4E6044CACD44657BCA9C855F65C1BC0C6460E21B49E5DBC38D74065A67649003679FE7472320C50A917B57A192B239BCE0AB9EDA5A03418F262BA83CF6CA11FFE237B8D50E74D93636187AE89CB8B7974289E8F3914DAE6A8719472E087BE859872F7050870DFD9D16628B99746FB03E9259CB3656B5150F1F696E5A6D7E66DDF1C2AA49AF39050D266C7DCF57F7E223375E21E620B05E025562E7BA892D65A9287EBA760D6DB540B43D2AA9163ACE5918E0B8B504B168900AEBE1DCD0F5FE50701E79D96E4DDEEE6D6CAEB380E13E1CF9009528D3E0097AC3857F6F6E90BC63C661D50BD1DB74B620395B10FBB07F2E715449DBC3A18E3C725681EE865C054EBA870A38F94A90B6DD02B6ABD82D85E9B9D1F9A7C3BED9083AAFEA87D5F720056D859B144EADE5188AB44A9DA18F16919C798E4792CB83FE8D66804779ECE4A83DC46987CBC0116AF423B55FF2E17CC6E9B828D63ABDDCD489A7F9DF63E77146A3B3F66548ADFE83A17A0548512CD8B4ABE524BED8E74D0FD53A4B951EF09E2CA1E22803E500B35042E8038EB88EACCBA5F00DB17203BB58114AD94978B444E8C36D2B654D3CBD84B8C9263F75E82C1E2EA6EF99684F4BB9394E31DA61DFF261DA1220A216B5ADC51F09B2341982D585BBD7D157C89D3FCDF47A90B4BBD28A997767776AA8B5603FCE50AAFB6BC0158C24AF22ECF07BFBD296772FB7CC788536433F11A62A44E137A383690D70DAB4689E48D4C29B10D84D47DB6C0FCB84F6DB88B7FD6FF3B89829300E84D09CA971FE87588CC083BBF0BF37EFDBD7F5C43B1091661547BC8E3E99F840BC97909C54227AD5147FD769A423A25BF6CD8A0B92B3327D441163725AC72E4D076BC52616CDE39FBA755E65830F69964774C3A46420B316ED78EB4EE2BA0A4E275484756DDB3C603CAC98FA1066F1F74FA08E04B4B130500DD7624A7D165534F1A560DBBCBBF8DBE90BB0D0764643D5A778DA5E72BECC1A0F93D98B09B866BA595C6CA93A741C62197FFD02307C50CB908587D03AE463FA5021B0EC122C1135586A5BB5CB66ABBB5C80F7268C203A5F19CE66080191522AF7E435103DF9DFB23256880903C843E70A8F84E170E49A093CA706EF21A4D77C75E3513464B3F625C48F083F6292326F714477F190A20913A4C2A00C7C65BE8F246F5879137190A45E1B8D9F168D9DADDAB5F6222956C2EF7F8856B9B1B5F9911BC9BAB54E03B4D4BBDD7A985D38C6A49BC21E7102BE9A7A70FA32733F7382536605B60094EC8B242C5B381C9085A8B2992AFEE51B220A7BFE87AB4977A0F521A8407F7F2D2B447E6A7D2C8E47AA0A7390D5DF10A098A00D9094259D92AF2298CDBD907D1227D29100F34F87A98C07D077ED0835F3FA858BEE86C16BDA9657D77A458BFFE7C4F81380B65D5DC29B8171BE012609689F9ADDB7F2CBE72583C3E00BD8BF8194D1639F80B8EA4B50CD48D54AEF3B46C75458C777E55E2E69B5C6829F69F3B381A708FC746F0C5CF214F5CE8FFE11E229058831F1B9B82A5A6F1AD6FAEE0B4487D771AEBFDCD03C6C1DAAA8346D4A9D51EEAE4F4276AF6B64FDBA4346FF73D98967AA351F0CFA3FDEE75C8AB8C6AF708E2B847CD32DE1287BE80C1CBAEC3864F6260245CAFDD07814777B15B047626E5C3BF5CBC19F1EE7B2B17D5C202CDFA0819611A845B35DFBFD41D32030E70A28D6F5688CF79547D371817175696B4545FBC1CC6075DB05811D273DF547A6A8942769DF375ADDCD52A0CDAD6C7834C71BF30382DDB0C433D35C46B1A758A8000D4570C96B88843A1C57BBBC915917147DF85963899825E251730ED7CD71E928701BB67293F0C6E5745934570389720E43418467C65CCAEF7213BFFA20CC477107B37710D26C9CA85508654CAF81A5B83B8A5C0CB0267D8C07F6F7F31E87C046F864BE38269C0415C63CA46E451801E38D893C374A637BBF1E4CF5C49083493CEB3CD4898427B9430E1BA771BC5C4ECC97224B448B8BFC1F7A85D30D4A4E8764B37F47B99621C9D977CDCA1407D8F1A1A4EEC4023CF5818A69D1ED81FE309AA5FABD21BCF3AD19306376DC23CE80967450461C49FDBA4DF490927360B76C2E998C22AFE3F796CD599D3080E832AE2193D839CF95802D5D14D4C4B640082789D48845074702CB6438031DF515C5AF987440CE4A79AF6C0D219DAC3647104664E010C48A27BAB12E14F0A180DA48F20C478817264450C37206AC2F2C0C5874CC6EFEC8D9719842E5FC7830CEE026605C344AA81D640B61A94A2E00A7EBB4FA961B9FE081871BCDAF801C69D3B71FC450C42DB8485CCBE3EF7448DB4D9F07F20DB228015B7D5A5E13C742996A65F12DB4B7DA0363625B56C04BC729EBFA4493FBEE36263D04EA3C5624E0407BC1529F9CFF75197909A075504FE6EAD9222EB3E7C17A6C920B9200586C0CBC8BDA23A7CE839B026A6971FFAB118438C35D6F7A9CE0B8DDA089FA4617A892745B0DC3043DD08ACE35B868F37D1F8B9B8D010D00E33794ECDBC78DCF1976C74C0699511C94F3D32D53913BE46EE342782652EAAFC71451C3AC775AF2021DB6696EDE8E006F9B7E1BB30A51F9B6FB93F38F9CE69E82629B9ECD3FE2CE611FFDD5B46A141B169E2B80F93AA4CCC130A0A90D9ADEA4771D874B975C1FB54AA32CD29EBAD3ECD8240CCA5851DEEAD86888AAF129AC4CB21C45624D9119708721719C34AFF0D43DE1CA7A7FDC0B27CC437753B2B3C63AD64451437A746739C946E26C30F7696A975546CBAF77BDDFB1864645709FE8774FB5F408CC45842AD9F1B59E6FADEE24649CA1608B1996ABBA1B529F3362119C59A6E444C922734924F061370C05EA30F42758402669B747856B774F2DFF0AA6B4E78B4B29CB43D6778A4123E11D078D81BB73A28D06B0B63111852BFBFFB151EB25E785286F418324D6D5F3F0E8B1A190E69DFFF713905D0754B7ADCDE6F8888BCF155B293472C18DA9E887D8AAAB068A07DF6F58D179C248358060730492E189D8FA20515A4F8410A81171628A06146A97964F1C29D27112E5738E7572FC43FE9D65BEF168B42C06C80958822821098B59A6E3622DB1B5BB79BEE6DB7672E277CD16D105E6B790A8DE2153040D391C628ED82CE12F7078411BD8B65BFE214FFAA946B68B5B9DE7C2789506EF60ACA6498869B3B5D0E57BF8C69C9E5FB6241CB800FD91F69FDD60281708D5E77835544018C543FFAA13CEC800E4A919F5C7591694B27E9A63BABA3DBF1E631C8D651737FDE4D2DD342A00E42934DE2BBEB6DE47E13A59E217ADE4E9C138D3870D6C1FE9B328177F80F934170495EF53022048B1504FFE23CE98301DD41B8E15EBB651962DF9957435452129AC4F40AB386E1DD59F4810C453E879630E56672AB53180AE8508013E4BF97213CEBFEE25D4C1EA04C48C5A771D73A77621E3C02B00A97DB25E3BEFDC7917BFFEF7B9237BDC9D3A8824C93B890446CBD9E8A75EBD0784084C59F2C0F231FF9A8EFF3D5DDD1996E3B44518884040E2FB7C9910D768D8F93DF5D74B9F36E137019F3BC744C2C5C46AAE6C720954DF41E7F70AA63F39D9AB95160027B4EA11DEE241CDBB1E719578FAFE4E30F3B6529D67A438BEC004055B7C332B190C07BC0DDB8117E5CA8076CBE679FA5B5CCA4B2AB30A5CB7927770381B68379996AB4F80D35DF38EEF23ED591A607FD928C86570BD300F941A1E44D4119AB1AEDC30684805E796F570F032A7C01706F2DC5F631D139DCB534A1B4C0D92B066238E6898CA92F38D2E4EF648E787C0EA8F07E479B73A3239C84E40816504E2A3A76F3E8956836D27CC2337AB191FCA502E449464735DE70942E2E697975A0A7103BEBD3A87C9C4BD16B552D45C6174F26ABC6570E076368A55EB7A08E67A9E720ECC8694BD7355A7C090CA97115FDA4A0F8E5F4ED160F240C48F0C52FCBACA21FB0F6CB1DFB313EE8DCF755A5A7329ECFED1A9D59055E008A3E8547A51A71AADE5C266C0FA2E1BEB7C7EDACA1D1AFD56F0DDF7C8D8ABF54BA8DD4941687E55665446D99760052D574C354753801EF7F01A38774B02CC6EB920569082B20096F3E5E4865C23DBD9337DB8715BB94E338420A0E02059FA15372CA66778DD05A20F016F63B4F000CEF329597AE9C17A3E8D3F0019111ED697AE6DD1EAE6D754EC36ABD5E898F85AF40D7A11A7AB084D8676CD886D621961DE6A5F2D003060B0C1D2CAEC6DF63DE38635451248CE409A5A41C9BD9A2FAD795F9CC79E165C05A8F11CA51E805EBC7FCBC5599D3CCAB64D0AF984C5FD82D683A7A7AFB2B09A730014BC253BACD6A1E236EC21E3DE338A2CF9FEC2C7CE2967447AF534F8D7A995B9EAD8D6108DBAD97853DD1756CCF7723B5581E8216B3A31749DA7C9859F60B27D63C23F04D959BCC097F870DC05C72E1FD77B64D5D7BCDF73C2592F0D05BADB5A53E8A1C4BA029AA71BB0C532F316BF9CB4DD1424E02C32700846C1C48FC5871BBE76AEB1A074890DE98BDB0B9C31481E666BA1FB02FBCE781A4C373E080F59BF93C022C05EFEC68E696111409F0ED11ABDE21A7F6DBE4434EEF78932C19997C5207191A9B2C73E4066D48B3B7DB6FF05D1DDBD371E7D2F339B9EEA1D3A176CE7AE49487833A8227CEBE36D90C7307DE4B9BEDFCBF26C66E8B219DD8D150CBA1C845F7E7278729C1064D41C8A956DCBD99D572473314A085605F9E08E8EA2B7C84B00CA3F4D4227CDCF3C8190BDF63243EC903624F14A6524C255C1BE992282CCC944DA37368263DD25CE639B3B664B19658DE30107CED3304C17526F009AF85B04CA97BF1B28C2505389A67F8EE6A57AC08583AFABE5F5C7ACAF0E1521A4AA66456682037A9E5CBDC0B36C05FA6D15C15BA0AFF8B5EA7743330536667F40BDD77EB51863644426C95B79B984E9818A85BDEFA436045867C4B333763A308FD959E1DBA61538DEB53491B03B8F50B2F20A2CE128E3D49850C6EC54C4CEADF410587E16F2E21AA40AF0379BFE759F576F109700AAC26F663BAA7E57D52189DF17200C9CE3145C8647ECB4A89B5DF79FE1884196640381E6DBED46CF5F2CA8653C9F1438BB30D0FD4BA26CB37B88CED895926F44D42BD2438070BB6445D5574D94E4AC7469AC33AA95E6D207E22876D174FD019A2E53D006D2EF2FA9058FB4EB80747066D81BF596D2A57BF4FF734DDCFAAD477E2CB5A24483C4B0CC4B67E3B06FB6D781A1C9016BFF48B6FF01B75C7C40315E3DC8026AB22E71D09E1AF8A417AB6F715B4A6BCBD8C64C7A8EB22CEFAE4282C05BD353072237F7F1AB95D3978306A74763C52A6F352C3A669AE6B190CBA3D88AFF57696EF559A8E7798714C44307A91951421DEA37D65FE0208A923FFB4737DFEBB0D8B6FE07D1B912388671939D0D0863C9EDE367EEB1F44FB7357827EBDF77F789F7CEC8A40BCC936DF8B63ECBEEF0BFE0D63E9A2C2ABA9322A56E9E83520875100749EF6853756F58698989FF0EB63D0DF84FFD18D2BBC4B20BFFC5DF59B135E8811F996ED89324A0126338FA8C0B10C6A9D21FAE71ADF3CF9497D04F438D1A23C3C5042FBD129A30DF29E81F7ECA5A28B74982D64BE80E3D5C27DD3AFFDDB88A3297C35E12CE373DF67C62012A986063CBFB8149C09E1947315E0B995D14D150C3E69BA3ECAB69D366AB7311D7CBCD17C5FBA7E79D4ADE02E8E4E7207F57C2A1E6EE3DEC8C2DE9B775BAC9E579E1DD486E8215D0E859B09550B4B33B488AA733D8AB9AEFC7BFE3E499DF059AEA8CF71EA7BEF177F0D904BAAAEF3684BACEBA0C8C775CBA46F71DE7C279E433A36C28736AD3ED7AC6F18219010C7F94FFBF983021BB68309F22353536580D84D898411D70EA41A692033D624CF37FC5007C7EF16E68D2A66E5D01E59F834E1040FAE78AA2AF823132036DFC8969187CC0376A24B94A748128F3B08D12A244D41AE00E5D5EB40BE4DA8269BF6E464C3A866ABB958EEB55EEE0B12D2A27EB43855F46E382460063CB80A204C62BA47BC567509CA2FC42FBDF60EDCD87A986DFCE4B88AFDCC2288B944910F73220DDDA5046047D86922B32B545A58FE845E587941F4C885E7753B7845DAE3886457A64FFFA5D740ACEA8B5938A6E5BD9EC909C30DB913283E558A2F2CCDE74B73CDCF72F1A9372169947E445DE59ECC9880444F30DD18554BF7AA76064D215F6F611930B1E3440490BBB714955FDD305A1997374B854BFA71434F6157D3DF58C58BD8DAB8519A5C067C953D36A6C9E3950AE9B63279096EAD9F1CF876230F5D6844EE278DC184CA20097290C4FEBE4AD67F7E681B13D2346D53EE9D299A8238367C94F8634039D8E476A3008EAC9E5691BBDCA1BD92CF0E14AE4586DB79B0A3C2E93A5CBE6050321EF4578D8A947A2867E13F8EEFF1DD8C91823785B6F824D1ACA20F798D0E770E0FBB2518A20AA0029283E65226008A18A20B7A2A76A2A354875AE4CCC3B0D48D36ED6AC608A62BFFF0A0FB1D93DEDA4A7EC066EEC408FAF9C6902D83F19F51EFFA8C7C4D7E409409F9286BC957B7FAB46D190EB4A8CDB3A79A2F034783E62E2BD879F1411D40B9C6F92848CD0AFA5A207773F4A60E101B25E41FF77629D84B43BBEF2E818AAD32C74BF533DFDF33FAE4C53C423056B47142124828E7CC5F073670DDBF465D4D12AE376F8DB66A089393CD10CA90F13C6F85F6A8DB1261AECB42DBD6D966FD41873905898619EED7F50E77B22A9FF459A68A48EBA523AAB917B61B36FE5BC185225E124D2343D289240179D262F0D3D5248B9A303ACDC0942B89286149B63221C4668F00BCEC688701CAA79AF7751F669DBA76524C5D9A8388B8521A38550C4F46892712BBF5000DA54FDFD3904AECEA16950049C32FEC543D53F1A52BF4C5AF06D74605B860E31FF6775FDF284D409CC913F985E64810A2815CDFAF4BAA9548560F315ADE01189F5F036D5EFAC4360015761701BD3D877E2BED56DA8F32C788D14E03673204EEADC3D05DBC82A8FB206052DC47B91E998780BC37822628EAE13BC6AC39A7DEE6E3243BD7CD6F2F08DC5F2BC5E49F1DE9F48EB82AA0C4B3F0B7EFAC34222E0D1F09EB479E7D893C1ED7A6F76E5EC497283C2E71932DAA7220CF907DBABB21B141E2E31817A5588E4A17F074CD9F335A9384B24B02147AFEBD9FA6888A05BE675ED42E49335E62E7D09CAD61A179D8BB090C6C6B4E6FFDD49DFFD2A214116B9720D544189E0F90622FA709100D439F327F04218CAD493ECBEBD91ECDF74A1CCE0B2AA0E31E508220C157B2E2A974FC2E9BB181D8D9848C752BB655CA11EDF719F97C3C068F584D88BB599AC5834CC3FFD7B190DE4758F95AA9F253D49B1A3BA7C17A155B888DB089DB76E80FFFD55033A98A3AF8D3C015B1CB8F5A08E84642C04F4D75AF8904FA1AEEA9C4D404A0E4274C7F37D376257514FC633FD489DA79D8240E073F74BB1D4C001DE15973A34F8F76F08FB179898766778015F37811DDC51CDDF377EA05FCF68F9A257E7757B21BC2F56F6B3D23DED9372C2F9E44BE6A9ED9137E8A135CEB7B8CE1561552DECFA1FDBF1C2A18FA4D523FD26447926E9ED003A0240F02F7153C7525B4C39B2443776399134117CF8268A9454846F4339D5BF70604E1F50486DC9ABAC58FB0A8B7D14F4BE4BD509FCF2DC29B9FD413D963E9E10332E46F33972A4B777F01D644555571148171894E41930F4C34E479C98110D8FE53931C70CCB05AC23570379E9D8B407E669137D254CC5448F9FE9E361BDA2CCBB20AC88A148C561CADC5BA82C668340FA3C5417E01DA39805EB863B774CF7EC0AFAD082F89860A973FE5155399F578FAC9F6CD66C6C5DFCBB1B04593ED190C90EF82EBDC3366879F291156B00A3F4F12508A8882F14233B523CC6605B046CFCB74CACE7DEBAF628E2DC48A5740EA23DC94F09612FD6EECE0C6D2FDAA6BA527850F9F8E682624991786EE56CFF2F1705A12A8B82EFE1B85E8F4DC51A1E57460ACF2D369E8F5FEB7CAA990D29FCD16975AFE270A80E613EB1CC4168E75A610558AB2B04F60804606EE1353B50EBE8035C260252CCCF99B5FB94BFED3D76E775E011BC8B45A28AAE8A1DE29BCB6A09956D05BFA6DF361AA821CC61137533DE8BE3B2491EDA3941F9542B21C49F6E5815F2705C7868F70CB130545B1341933914B63DD1374243D63287714252782BAE74352AF95537048298F748B269F6C990269B04F549FAD3DC1951F3694BA896F8814CAB13553222B73DEF61CE432F198003A3E67E72C0CA71CFB2166234F14FB7B3E7D992BD73C36C0EF810273EBA4161A8F04D04E5EA9F115A39E575DDFE7381799C8A21C56777C06A85B063A2D11765836CC054C6F2C39BA12001037BC02EF89957A74DEC9233619CDA2A8EEEDC263983D1B12C32B9DF54BA4F658B196116DA68D02EB35DC16734976F3EC69F0B1DA041F519E33916130FC37D5C9875BA3C5E03F979E24C7DF33DEDD154FB6FAF1692D1CFCD1E0499CBC869B441736DBDC6189048CD3CD2EBB4C056F65C1CDEDEBF00E0070F6854F4D780344639F666549AF1C7938E62B2A1E1AF9F89624F9FA06C89249CDF782FC303232F45C3DCAF10011A7B13E9D78C02EB100BEF78715689C34E597950A52B703C978802F464F0A55E949DD783D03D8E207B336902DD1801BFBF85D5DAD491E32560220D482425C85E309BDC7C78AF548350222FC7DFC734F13A52767169135F2C45E0B387ACC5195E7EA0F3D4033B8BBE5F6CBDAFA38A77E71F4A7E245C88CFD0374398CD6017A025873794B7D85BF14A4765859D7910486A471E219E7F436EB5CEEEA96CB783EB11CD61924F8E2C1C5C55271E51F141D8A59AFC774B62C2304EF715230B18C30AD39D213E0ADA2DD4BFB67E49185BA27A201244B01F0E0F147EEF8B139A200BCDA17C9A9A053A5D864080F726ABB1037DD93D5A7584567D9EE9618E90118D20CF03B0C148FA4C276CD7F9C8C82AAAB7E355A92C96792580C1B0E1713FFA3FDA576FF7C90DAF34CF29845F3FFC54BA5200C9B42CD501C358DBDF1D1F9D47375DCB0EA4C0906792D82F08A11D138A4BB9BAF536C1391062DDB1B12A41B7B16D48B0FFDA59ED4519E486A51B2D86D43AE92C63DD4B0DB6E5F6EAA6A7363C01DE87EA95CFAFFD378557F085AC1ECC5E6EE1A917111C92BD57603A9FD40030B9E0E4A66B49DCFF49E3A648CC3130DF95337E9D1611B6F131FC5682DAF6ADACF944ED5C86350537D3703BFE9920C204BB8DBF04B976B01C61058C3D376FE7A2FFD44627CB6B1D8390B46111869D48C95D1FE90AE597384F02228F737776F1EC65432FBD82E3DA43ECE891E83BBE172ECE2DACDDA3C029B9E5F6DB1A6E20422B2EC699F54ECD2AFCEFA527F5E22D739430C8972B0F85253E72A8074081CB4FADFE73DA19ABEC63946ECF3B4B3CE4332A3666C4B23A7E04DE8AE2703A9F90B7B4D607AF08BC741E0946CECA731D0D1356145FD1D4E695881E557457D8B7750FC889829D0ABDE5A20C2BE4D4EDE29EAABEFEED491501FB55F9D23FF0244E099F456A494C2FCD7FF745892D7DB6D2BFE53C68F974B2A3D101906C5C83CD58A7199146E3A16C8C3A12E00A12135AF3B6671DDF365C3A2D1DBEFE744FEDCF33DE152EF4AE5D76DF094D69B9AF1890E5840F2B7219D35447A2435D3D62ABDB6ED2817990AD0ECF9C74787FC6CDB56CF53D9D7FFC84A46E6B098F183A2E5502BE257D740792AB40925247DB4CF0EC31D5235275519766C6DD210A615E413C2A00C4DCC0CED99D749274E1AF031AC06B5D41100818016988DBF08A7531A90B59325B4CA95BFA748DBA672037EB6250A832C7552FB0241194529226FECDA5006C33EF33F76D53FE95229359CF70BD983A07FAB71A94F7C2F6FAE25D6D9EB2598E9846FFDCF7EFC667B409762E3814E76166180BCD3899C584E4EAE20CF944C06C127F9E8081ED72FEF481771191879FD40F77FE041BF166B819A879657CF6ECEE1C0BE6ADA51B6A0F2618C1EA84FC0494E8D25E9B90456D187418206E8AA93F8D703FB94B6B6198578323DD19FF691B513E30204DDFF07B9139249C5E91DE5C5110BC39568CEDFD86C015FB65BBFE9076E5AB998782C61F60E48A4D7C317E83D6B65F1A7041C0368412C63E8734A5616968C5323DEE2210B5AFCA24B84BF6FCE8721419A21876B1DD58726FDBFFC7372985A412E3FFD4D42A3CB8B409C3C8A89A0A654431DB54F68B3CFBD49253567890C2D6EF2C9151E55297E85B1541675A16312734DE1240302D9139F628174622DECB851EF92B5D44297E981F79C8F1506A78703B4B71FF66C42A833A9578DF83A420D83EAFB7E90E6E4F2CE76A8995801F27D8BDB957C721A3DE3B8FC04172ECF6202B77699094B023026A196EB1745BAF9B006B67435FBAB540D5AA46CB1DE630CE1226F01374BD237F707E854668092D6992430D3604522F1072AF0A223B33DE21F87CACBF4FB2C5AE28E1318125DF2A44096902BF38621576CC03950A601737E4A091E4EA5CA7FC7C4169C7E33810C16DA0A00000B830CB09E2C8472AB0801835355C5CE9157030A3456C091A18FF896B2E4B7464B31247D14185588306367F3131BEAF7E2A697A042C516C6F8223CE897983F31FF9A3C48B357E4D1EE445F9CB66962374B9D71E4344A6DA9FB8505A9D6CFA91C90AEFF66D9FD6D549A78704B19663D33F57ABCD9BB235013C3045145FDF28AD282D048537B3E6E764E710C65EEF8197CA2C4CAAA578EC3E0D10A62676402A9F20A73C53A660EAB361D64256BA5D69A4320A1376DD78D132B68D99814529979B975DFB7F21F699D04BFAB3BE78AC72C47D556B387173F4854E19CF0DF9BF6F5B5426EF59E5A8FA5746BCE32CF00A67D1DC0BF173AF3E2BCE4959C0D7FEB5367B42BE366CD7AADCEE292E4544F5E81BDB78CFFEF93EDAB862092B3F127383C2D594D9A85D15D1DCB17991E997C89BE8E3CDA01A879B21376FBC224B2C1DBC088940DEC95F9837A40AF69C7CE8AE446752A1422906E25A8D20AFC8BF5FC4DD753C23D543F238B8AA952598A40CCB9C3355DBFC6B0BC0EC3092CC7EFB62AA2447F9B542A6A281D5016556866BF546680E05C443015BDB9D96DBA59A38BF112F75ABD4BE2D3CE9A1AD7914017BEA55B74550EFD9440903859CD92711C9D08B28071641AB42E49329182DB358FEC56815D659527825E40E5905D4843A53627FC94E46F716C1B2696BC1FF9F2E9667BA38376295AE6F61261C3402BDF241B71C803B3A5F47257C7FE436E4D005F3A26778A6DB1306C60E781F54950C6CB322E8E4D45608F87CDFAA6998E6E62686A05338682CF0493A1397FA2E16C185DD4A341F6B38013A291F04DA226D799A93706EA8BC4974330C2D796E4AB51E51261B7354F7BA18B9C6838CB1A09A99CD5AB5D6366B3AD8615123C72C0CF9171C45F49F553E0F3C1D67739CFA321D16DD74A871390AFDB13CF7A901E442994AB8C7F2B1F47C23CFED3D84F3C24411BA1056133157A55CFC159380D3826045BA39D26C90C515EDE1379C34C27FD9C9990AC2A3545D8DD00C313FABFAF52F0CBFCA848B7D9A849A4B860666206EDAAD22CC4136839DF430856214C07ABDB5FF5A38C6141990B6AE86E47E6748F30D92D9E007C71E5BD5CE308687DCC57226233B0635A76E4768D5CBCCA21A35D68ABE55F44F8A00AD281DAD5512B50C90D1D4371A792966C8AB839629BDB0764ED068365FAC21147E90F535C20D1C51CEA088ED498CB4E0018212AB18169EB144128FA0A60DD0DEEF88E56A146B3157A4C2273BE4844A58FA3EA7C2ED116B6700FE332EAD56B016298E79CA8E46B24E91E19862733C9566CFAFF01A72241B3645B8FF0AF169888693C6E1A111EF44163FC23828D9D11522E8F98901D845F6150679E21AC29379C8E1BA913B7050B777AC04545EEDBBC24B387DD02AA8B7219AD2CBFF3DDB2780A0F446547D7792D8E50BA4CD6B00D3AE3D7C939EF6F47FB1A7210A176A77B80FDA54BBBAC60B487097292205C47E425EC489AD8961368BC320E5D09E656AFA77996C50E8D0AEE864B7D93D282FAB17B86CBCC5691A1625375924B632F33AB514347C78C80B79A3DB67EE04D16BCF1461BECB195F68587130A6AD651392BD1E5D22D857512AE9E8D309B372BA841D47874D290014C068D372E1A3CDC9FE90D5379E37E95AC21E205AC4FD4219BC857C13DDE5371D10D994FB3FEB620BBB039C6640034CE32455DFC8A14DB058710268D951962A4D3E7AE98A6D578CF57611EAE96CCAA7DDDD0B1854ECE3B515FCA6092DD52A5E2AF51AE3D3E340DD7A75C767601F710605BF279D7417B03F4AA9D8CCFA3C729D4D068B5509872EFE895F30172588A9084CA68518B9FD428178D21363679F6ACC79A35F1A86ACF56DEBBCCF9C3BDB81FB6CFDB9B57358C41CCF425D733A38B529213CE04703C0E48B1C05E3AF5523372A9509AF9E66441F2BD3E6D3C8895F8D749EC07D0E7BD644ADC8582965E7D2DE68A7580E8DDF3FFE602411FD8474C9A3D57D7E8361F5488C0EB98586C5E04E7161B46AC494D9D3F605228D985D6DDCB44DDDD5AA2597C48853DA5EDF77FC196E3616BA1624C1A822EFAFEB473CCEFE1BA9E6DFD246203E32C0C12AA77C7E2CC3CCFDC7662F06E36329872029FB4EF28A1B7073D978A8A2C4A5121E391CAB9EA549F8DDCCFC73B407037435513ECDC7107B7C31739AF90FB95AE82936EFEB57EB9ED36B50F76D8FC0F5E9C14BA4033677702174045B1A8EFB898695E24ACB92E070DDF170E340045614F2B26AB172242462C20453BC8FF4A1C0D67AF0F6FBA710805E7427218BED1AB198078985404A07EE1AD8F18286C5AE2A5E68143B40F1EF91F832724824408EC9600366F844771C88F1AB9850C77A295BB6089DFF702E65D94982DE108A1094893E465A1EE2D2A0247E9C1D2B1E0619DBCF8E8CDE19761D60F16574BABBB9BFC9004695054BB0538E4E5B2231C77FA45128385E5A549994E2565E45178FAD5B3F498C96CD42D8062FC945BC2F491ADD070394FD4B2C10038668A06DD83B0906FE6B9DC0149296279E1D3D37941D1C05C0338C8C9187FFC10E8C74D4C0E5A5438B44A35BCBCDAF2C688D1DC8AB226E2A7A9A0AE2AB1048091BCA9EDBE5A4328C9497F56CBE3FE8623966F7C64DD4B7E18B56C23CCBAC6BE4C0FAFEA953B953C6F6114EBFF9472D4B216E9FF813F5604334EBAEC9E6B583FA23E3B17D4248385C8415CFA5DE3107F8C2156246EE30E8852D9222107153F5D5B0AB0123FBDA39084DE1B002685B96ED3E899918CEBCF45C92E2946219C2BCFA63640CC23FFBEDBF32744999C0D26758C2C9651D07AC413E1AA99AE2D9A940AFD95F22FF7CC8751DF23FE61484AFF3F322949AF7EA1B0A3F49CD8F73AA14BDB9BE44C450459A82D305C8577401AE8C35E1FFA94C4F67C81BB9D06C350508C6AE2A9C4570CDBDBC97822487460E5C3A156B4356396B95BEC59E59CDB1796B3CD6978BA1C106A5AE352C3730856D1C78ABC6D94EBB3D8C691BCD232C293872F780B69279328687BAC7E09E351D5B844CEB9AA81E9060C642C27BECF48B82D99EF509030E0F0719D09B1BAFCEC55269604B8182A504DE63DBBA6475DEDEED1826B05E0962FED3C89C15C7C1749FBE333BC8543374FAA4F52D1ADA867BB565F2CD0292921BB97FB7AF211FEB66EE9391EA99B1F857D8E8F76AE6BFCB494161BB177DDCC1D72EFE1AFC77A0DCACC0D8745C54F81233F6208EB292B23BED7E7BF046A71CCAAF96DEC5F6039B8C44AC256BF3BCC2BB491D9730F34838AD83AEC5D85DAD1AE6C42490976CF2F0B50EC53CB2C75D673C7CBD53E44223D0EFAD00E34D1060ABB84D477A2349B208831251B0ED3022331F4AF9208A13BAD5F71BF91F8AC970F5C2A404464EE2F1F3E938F923562D49C216A3611A761A5F7B864E56582C26883CD62C82A8F6191E69340F4CFFE42642A0271A19FAF98650A8A892EBE5D083CF8AED4E58E285CE7539B8DA539C023C1233E8A3C742126279006256795F396CAC82F4D05B55F08037D9BA73C0F5A37DC9C634C757C1A078FA25C3E896435E9A2CEB1F31F9FEFBCEF96DBCF3689AAD1C9471B988D7EB929938549EC1203D44478A95C2E72D235D9961004C8051FA46BEF2EF75FF880DD8980F5F67A9C8E1FC74B9DE20F7030300ADAC65A5EBEA7D5F1B1E84239ECA89E391A2B51637183ED7F1793F7C1EEED3354677C457A97BBD2624F9A261AEE987A6366275E9F72EC95BAD86CAED0380449A0CECA8A0A43CCECE60291208A1096F80DF94322FD974464BBFF12237B27AD84C2366AB49D28C3ECA5BE298728523942475235CDA7F74711BA5C4B70B4C8C9113320E150AC7A6DB838F84770AFDB0405A45742FFA91547DFD7B1D5B3A6DF8B5F6510D2957BF79903F62CB6DD8732664FCD30B8BFFF07B1E6389D20626D64D50864DBB36A89BAA599F02A9D7F019D4496ECBD0855E09F7C141F2B72DDA5DA01DB1CF3E3E232600F0D29CFF7EBE2500B03F2513DF959FE5CE41F0CDE8F6D48F139922707D71B4A50D947CEEB25C84D296300BECCD1D4506295D8F70AC31D39C600086D5345E0DF526DCADD38CD0E6C9F50CC8B4B69EEBCDF976084994D1E39A18E9B2216B84EB1AA3B0AAA261F2B8735828ED02F9346A408D8B41286CBCC3D34B0132B40068FE9C60F6BE2FDB61ADC360BD9A8B62AF4CE40084018111203CFC20CF32E220609F6CA9E966445F2D46021BCEED20E58A70DD791DB46375ECFEBE3AA9E10C611A0F2681229350A40B367EBD71D34625B70E1317EFBD21AD0C13C1A1AC63D6B5726218BB88215D1389230A697B8E9433FD5ACB97DD8B8E999A6189BFA5CEAB0843E184DA5F71A8ACE9B898D3C5333C969FE0718D9C288D12004FCB7A4371AB3FCBE496AC46E4E937BD5822A97F7FB28D9C4888B0AC8A09F2363969696E80130A9F1E2DF4199259F52D38BD601C4790000C139EFDF6C6167A37EC628F08D06F1AB497DB46726911F6551F7342C7E3CEE8D8EB06080B65584E9216EFF62D0BEE14E108054253B70A4C5C71D47ED9407F6241A9410EA3174B7994C4C670E5C315AB072620952621F573EC2B961157971768E65B19285B48DBDBEEAC48F596FFE8678DE8ADC4073392C9A6244A1A1B07FB1F88CA9497DFCB1212D48ECCC231FC7BA9987A778B878E2E64DF0409E3E39E013FD00070E34F80966F57351F46ECC75D682D06575523B3AF5A135A5D9C0BB0C72E8B9104740BAA1F4B2C67AAC6D39A5190FDF21E872F645A4B13377705C7029256BB36EF5219885B208300CA6DFB4D9BDA5B66984F905E6B938731B1F12570F51265BCF279BECCD60F4DE4C01D30F38B5F978C5E12375307203C4121C267400F34920FD60BD551DCA52FF5DF5F48962926DF9B58172406EF459D5C2FFD30BBAD2A544798CCD0FB2B44B44991C75DA0FF2C60188506575C918EDEC3E45ABDFEA504FB8AAF4669385E9DC8BA412AA981330EF90AE1FB6DE45B7C91D301FBB5BE31041243579372343751E3CBF63A9B803A125251111446EFE2FBBA4C2B3255226634B41B72590AF61BDD2A9A30DA635DE20A018F411CD7FBCC638C117B52E17F128495A390B4E3B097BBEFF0D148FAEB82CA1E630F534D9C868A462F189CF63230A12AE1661DE95CA1D78FD3354BF584900F72AB61144375B1DF94142695B50512AFC9FCAD498032284C306D28451368979AF734CAB269684DC308E65EFAB8F878F66E9918721BBF5709566E393E59F95C7465364C68D73ADE0CD6ED8879ACE938E8BAE7DA545273A514B744B9DA5ED840F49F863B9C38A5FE8F1E1FC30AFD8C9F6856535A292DBD97F4D8EBDAB6468AE921E4B3BAB2C0B869DC7DB7408164F83F604533BA262E5A4B2857EA46776958A491B531F0FBFD5335AC6E44CC8C395B691CE854396C4B3A2A74B469DD17F5E6B59CCC61BD927335FA1C6A3B1854F74658D4328C9C2C011DDB988257453474E40E3778B83A0D6AB9B9947746BB0D82E45E673C81CD20DFC78A9885E8DDB9751FE583ACEFFFE500EDE69D086195198BC6CBD9C63E759EB38A87B8BDF0283D4FF4B6BE3AC94F00900F5377D6B66C3E886533E776B9F2BB43566BBB2CB4CFD2997284118D8B3032C34840098C70624AA44E08301EC739882CF1442324A0470CB997830C87C95BF8F5A391EB8EB13D962927F2FBA2EAB407F6AC77E195627E2000E8360053029625EFB9992D4EB259459F22944ABE2CAD3BA9737957CD574CE64494F945EF348E25F373C22E2A6C71F5A9875E8EFF0938E3405AC3A9601799B2C0DAA37365918D4CF8B03551360EB92B9799CC5EF439414793586FF966FE0180A2224E1F4D3DDCDC62D68FCB3D48DCB8447CB25E627C0CE07DEC66824BABED1B6C43FB1718DFB67B7693EDF6A6B3C4B864E00F65B131C59C42E42A87FCE2F2D3DD60102233550A87CEC579C9EEEACC386479A40AFA02DC01C467096FE3E7AE647F7990458E92E732D7FB0F29327102C215716D2185D23D56D5A305C293ECDB7441931602DA8B6277E9BF9B419295624E03931045669189F38B8071162346275F00856AC3ED0C9B76A4D79FCF0244B0DE0AA97964C18EDBA6A733CDF7DFAA4262022A17934EEDF2FE973BA14FF4D4C6D8776A1D38C27833BEB0731B0AD0B167DE31CA5C9521238BE3B545F8E7722B426ECF974C48A036BFA89FB6F6107CCA9E273E51EB5DAAF9858E31F052A83C0005A2188958FBE3C820EFF237DDD63B98F400E912FAE81D0748444F10C837402ED60F37E60B549BB2E973B6EDB97272440D765AF16C4174BCCF5E885BA5584162342730AD609B7FAC933371D3C5DCC639D9ECAFD84E573384158F5B3C7B8C311F468FBD2F24552B6D5EE496A37A2ED7A6A043659A7A604E5B6ACD8B04C5160C4D2C761A252000FDBA58991A4BC73388E864C5EC11E0A088F4A55A65108F1E298BE1FBAD3BDE136B182096C319EDF9CEB81718167BE0186987CCCDD94776F5C0866EC67666D83EF99DE8E26E681364225A02A09C5942F91E0936B46EB2D0B2126E3A08BCBB390881B694DA9644E1270A92020BD1E43DB6D420FF4A402294161E0F160C4BBA5552E33472D33A3362477E4EEB22A609D2CFAEFB39324A25A87D4EAD18FC133801D6B08D81ED85B391732724FB7754342F0982E875288385D298B6CE6FC4D9FA86D585AF20E283F57F7CD4A55A0CB52F566B1226994F44EA96C9664CC2DBE1838D47AF3122710BBE35F8A2301DD30E7D22636C8B10CFC1FC688A3E6C69E38AF8BF81076E424B79BBF028B0F5E38EE3DA5495DF9E25C2101927F6E15557ABC6C8A26E21EE6F4EF25619DCB13832EF7CC7DBFD3B4AAD5BDE10A104F805080745A28B9506842C482E1A92F75C1A9C3751BC0DAB432B1DFDCA8EE92D70D65B643959BFC29358611B81D7D2280306161381CAC241DCBE2DEB30D20BED1B78924E163F2654857FEE4314D6D24D81C2D9CC9301DEDC39EDD62D5F704B708D2BED2CEF13C73ACF280B21EABF0B3B679582DF9E294BA383A00F622FF5310E83BA9E5C3F90201DEE25F33F36FF7EBCDDC141319CAE56F9B0EADCA925EBD4DC6153394F061E03F17426E6CAC171D20A3824BFCC9A9A9FF8878DDC6C25F35F4501037E50741B06D56877F46E8EADBC1CE553B60B1781065DA7185AA447C70EC4ECE89B21FA286DB0B6F1FB1A2B0C1E1D674D0AF3EDB6831BD2799C87121766F7BD8465D4B5380418BD1BD4F4B096781CD914FCA4B0FE216D2789A1DD411299B40F7765744978611F024EC10EFE4695986123414C3DA35810C47FA9B8E635B74A1EBC58E1DE8A240F07D2B525AA99760392D172B9956504F676F6304BA9DA1F261A969C3E380E3310AE0B872D4F6E1C5EEC6363D5F681B5FF5C4F41C3B3ACF594FB29EE4FF8883B9F061A2A1C2CAA8372F9EF28093AC00429F6414EDC283A52A88761DEF33D1B35A6FDCB72F9BCEF7828F4C5B73B363F5456BC1EE115F4967AED61CB769237F99E48B78B19F7B4DA7BC7C82E99DDA5BA86F08F8C1798D609B0F1E47F7C8F5B4073092C5E964382DC52FCC31FC1BC39B796E3C86C1B32B4C2EEBAA5298F8C3B3981342347AFE70302FBE2A929D02F95E8CAB360C3DB6A9EC8A13223428B0D5DF0130677C92C5E3BDB2B7CDE694658E1F66C3CD757059AB989358D57A6978689FB3A5A2A815BE055F07A4C740253502F9ECB6630150EBEC4569ED6C872677862797B122F42AC8450D39023A32C7ABAE43FA2E1005CDB99550917CF942587A52CCF40110AD3E9C31D20EA67D7328155C5914BE633616DD122F77A8C146F00B8D20EBCA9998F548AFA33A4F78DAEC259986F25B45D406BBE3B68243DEC4A9D5603D96AC8B6C707C9B0BEDC6FE5629B53CE0F5B7E95C6C1E0C98B51EB0BA6D3700DD8D8A5812BF125FFB524A24B84362CEA826A8F6308561033899974C112A3FB429A953C8B0616547EF2AAD908B8E3FB7B1A0B4D0082ED72E419C67F501211C861154F2AA02A4E637D76572762BA3FCA851CB5EE556EF0A530434CB6B2BED11D6A04C5FCCD1263DB0BB6AD328740E5992518EBAB6058FB79CCDC00167DDCF23670EC3277F4EB60D3BC4A33EDAA2A6194940CEEB475E57536A01C7DAAD06180403C441BA514E2D2B9A557E62FE7A6FDA79FF0D4317B9729B7F269F018E03557D6E90C4F18CEFE7A748D8E62BCDDB4F9DCE86E34ED32084B880314C3307C4EA4418B1F5B0550C598F4F41CEE7C3815BA00F0167A5EDFFA3F366D0F452902A02563E4D3AFA3DADF9A7BC5E7EE42E67BD0E5BF87D2A39BE72B1C296CB3483C8FAD6CFD749DFE4A8BB297ACFFDEA01CD36B853EB3B1BADEE5EBB6A2B440ACB7FF9E66E7EC06E5A212F1748C3AB9CF1F974B30F8F6D6456229632068C0BE1182E86F5C40991AC4985170225FCD320FE2E4FF6D46825A2AD839EC25A3C51E358CAE77CDC4E0B0225853BC7D39B1C9D89188C8BE2D9E1751B516203B691B82C1B8B6C6F332CCA3286AD612F733AA5E4131ED976D8D8BB63A138A992A4D3232CB5DA3717D1AD93F9153B84AB8114FE96E92A0E14CA1BB9D482880B1A2771A7FC51D6FFC0331CB22322669AF952DE3E1A5ACDF694CC700C411E5F6257135EDA931F5C5E9AADC3FE78618D833D97999C24454397E2268346AAE28BB8BF2C604C284CBC71F418C7D49A9A6D6BEB5BC157077551B3B1F3136EC5F0FB6E98DA63EC0175A8AA40F8D48B34FB2FDDF57A8C0E87DBE314787F18872F8CB61D1069987E1032F9D3E99740B07108EEB9BC46AE9ED3C8E5DF6421FA91E654BDF6EEB4F6718D6C2316BAE19CADDCF8A198D5B1DA022232DF64F75FB36DE1D780BA71DF1F73562275F7481715426B942652D902FF9C33B81193FE044DBE771445D44BDA7CF29DB7F68872399B91BE8B2A9049254587D3C10BC0178548CE0B0F0CE772F9FAB17E2AE3A0535B6438EA4D7B54ACE8D5E94A63E829B0400BF287D40008D105AB1A65ADEBE0A5B37E78D3882F4765C96A84EC5FEB96A7D155BE0DEBCE1B274B49E8138F66D36E73D4D528193BEBCBBBBC96AC440452B25E4404F0E35E16BBB26DA2D7612144632454CE9B46274B55083AA5F2EDBBB4EE36644EB42D7D1E8FE3F2EF1720DBA7E299CA5FB8957DA1EBBFEBCCECC474B08B3957A609CAA832EC85873671ABB326A24F4416B13CBB4791B5CE65729FDA64DF607031640035CD592BD3A6F3318A50803CFFA0B7571AAE1599074A5285C93A8C146806F3C3B27594BF99FE50CE78317D43B37793002E25104CCF5957845C357BEC9BC43088D2DBC18D86AA84EF002449875E6FCECB2AB01EB9B89AD06689A096A10E30668C04B31135E639D934290EB33A99015CB88049C1086C68771A09193AE337EFDB55784476168D0C961CC0B2CA4BBF0D16F7B21E3186CA3EA7BC078790F0034E4E8014913DD5F781F66CEA09D1FDEDA3539450A2C419FD57BF033F8B2C75F694D0EE2C79D0BC1696C61CF2234120291410C5916FCBA5E330357B43FA40EF7F5535A707C7D3AE8D2965D6424B973069F12841DA265CC739082117FB6215134711D607E89EA6197A101AFAB934D8B27A699BA3F526C36EBA5C86AB479CBA0AE565D8DCEAA283F7F5A62AA06B5F003D9AFA38B4BEEE529817418D29402A3B3DE15D863788BDA2C2EAA824DD8BA98766CACE49B90E28D370B7C7162150DCE9AD7945F04A9FCFBF8E0A434F314D2BAAC7959DD9561B135EB8CBC6C86C1CB4185C669C5D9F984A142B7080CF625DCDCCEA973AC8995BCF9D371CE7A9A8A034BBAEEFD2DAB86BA0E78E882E5852561F0F503902BC12628F6C1ABCD152E671184BF923200CE2D79DD9129782C23A23280CE053EA58FAD903775F4F9AC84C6647B0A58F85C28159683CAD0185B702F0B075416FBB541E67787A045DAF724C669F0E738900E65E3CD027A2C97B41270AB1C2E629BE1FD765FF4688D51C9FA537F93785B856DFD2109DDE628A8FC4917B7F01B7E450D534C3A54FA6652AB40731D8423BCAAEB1DABF796AA763AA72BB1CCE6682A247E0B201783CE2562787D2F9E44A2F633785E27DE3F4DB3BB50518A19E6977D27BABC10C02599FE0BCCF5E7C0C5B888AA71503E7AB8B08200FC0D994A5DF53FAC562AAF1139E5A566B4EA33B70DCEC7A1DB382B971A90FDCB0C799FD7ACDB7647C870093398F3382F66A06E9D3FDFDF81B4374A1BD554C6F013D2C82453D2EC3A7D5ADD0A1B39FF7AF116C5A817DFCB8D40A56DC1F53C523ADBD98BF21B95488E614349FAE280C5AB41DBC58752332B776718D2D00E203A312034B72A8E6154E9818721BB65B107280BB574DCC655A74B8EA92D512C1A78DCE67F2CD1166449530B98D43CA2A1F59CAC641708B8E73D4B67A399780CA910667A0D656FAA838B276E9ECB6620488A3D763A843AF99714F92B92204B0C7E6725B6E24DF84EBF84B14BA0DB8B3BC7FCDCBBAC4AE2B42A77218C922906D79796315F4E1F504F985038604CA3F4E512B39755F8A0374B1F3E7EBD8002B71227FD8559310D43FB7E424D50F551761120F9D6EE759F587FB7B335D73F0D2FA81CD90539390E6DB7881C199FA849B86D57F4F61D4E9A39D923708136280193CDD73228C350388F80792BE0AA7016B038D238AF055BBA04AE35CC0CA7241D82306A873A423CD10E4A13DC1D099F525033CC8682AF4002472ABBA73A546BA1017697768C52A77981BB39B193F2381D2DDB6FDB170ACA4AB6BD6C5A424E542C6C66CAA395CF7D225A2CB3DC7CB4911597444B99322FF4E4D664228B35C743B8152580CF0FEBCFBAAD89826664EB6D714D1595137FFA26010BF090AB7A2C40B3A1FFF538F0CCFD2F67E817624F389358D72A2C3DDDB81A4A77A9119790D4F2EA0E20811C9DBCBD138D41811A3119D6E8CDDCCD8B3F4DFB26C4108012146E17D9A33E26CE54F1AFAB7D0E21E11EA6A34E80277BB5AC604F1679A1FCD66B44F3D31214DDBA38A28D5517A1EE098DB848AEDB4200D5881AEA47E403A78B799F9A260B3AE5AAD17EDE80CA3B4B64DEEF8B994BDDB8C38F51A33C3C690FE88794CF56C2D3B2B362421DB80ABCCD594B5015575BA533AFF159DC9D95B2F06B4AFD1ED7DFC5EB4283AF716D2173FED1E111A7F9AF723ECE8522A3075452864E740AA91B7132BC61E772774B0E974F023C9A13792006204B705090463FAE00EE4266ADE677DBC0BE5A978DC91A65F3273E75C9DE8810C3A86FB300DF473E962FD5025B800143CE28CD5A64CEFA1A7C536800E36DC0033B5840B62F444D3F7935C6D0AD2E4C00015D73B51C70817A36CA6B1B5355A499BB3054C9B151A52F8A71ED65A5A0800FBAFE2637691527FB51B51F1FA0920DFB376ACDB74FFF9554431C25C496F27C8142DF92DD3BC3EDD3AB327C984F94697DC8301E540A5F9D36B94B903787ABAA611150EF23F635372B4F48E6B5AA0AD254FD9A313B1316B8F704B8423688DBDC78799FA0AD2BA42F7975C8502B66DF4DFB5B11C0EF58504E79142BF6C2BEF4C012942ED14FD435A26B2ABB6C9B15589AE1C8C17C382017A2C5A9BC15477EB7F8FC6E332560E46C80EC3B47D8CB93A6E563E340226CD62C277CB3A35F2CC609609DD7568E1FE7B82A6654AE4FF5524EF16F30FB34C006EA1EF93F500A4D46D91B826B11961DA65344A3C9E079565795BE36697C944978E416350F87B29195FF24CE28DF4311FD8029CE71576F571FBFC0182F3109D727ECD0017E45E1FD738DC2AB242DA623E8DAB59983BCA5F47E0F4356F97274DF284C03344AF1DB939391E56C27EC0A31F1CBD11828BABB877B628326F970CC2E62BF64828F84A44B4582FE633AE7FC83550C3553E9136BC7BED69D995CFBEE99D9D9323E59844AF3EDCFC3DAC9EE9B9D69F3E43D612EBDB556F4A5D613FCFA3701F9974784F8B1347291875C81EE520651C4DAB7F114D588764222CCCAE312C98B39F21B140D3C720FFD7A041BF2F5158999529CC291258D222746EFE7BDEB69383CBEF97085308B5F1A3C2125D6A64BBA7AFC767BF25118FF0727B3A91E8E9A2C89D3FAFD35FBC771D8326911DB16DA9ABBC87654AFF41FEFD471ED289A68F8A551DB5ED1831EAEB1CCC9761F56A0B5422E9EA69276BC4D69EFD19293CE53EDD9BB6B4E2280256F31FD9139B888D9C78F17C149CEC7C1792C389E635BB04F97BAECB30BA11070137008DE630FC1CF248CC05D9CA12E34C564B8F50449FEBDCB02D2254FBAED4AC33AB1BF577B41423B5803876B48B8A1F11E7C82D9B009820D6FA35258865CF479B59AE32E1A104F5EF1B0FE48AE5863B9EA5237DEBA79DB714EBB1A26B46D75F1DCC4B29A452003DC3D46638EB0A99062A72067E1999E25D77F71E28028845514E94C66AF4FC0180A369A74091DCDD47F790978BA44A600953BF508E6CB769526997A510212E1D1B9CBD5367CCF5EFC77626132147613AD8BB16C42C161D01B045F42CF0F9C008C5ECEB6EDDDE412FFDA4BA5ACA9ACCF42DAADDF8AED793EC20702D3D43277D5DC8F3FAA3B395D29B7735246B6E6995D421C69D3F0A22314AD45069F0015410B8DC4C41D4C2B980F3C898AF425B52DD16D1D890AC83B963C5D5B36700483888A07C0206C094A996155CC3BCABCFC9DE19F9048933D967283E4523B420F04856A8BC8DC2D3804EB4D95F360EB50BF2E73A8ECD4974874FB05197E1B41E0C3F01CD0BFF54BE6AB6A9AC3E456497B422078F779B82C4CD1A067ED0D6B9568A68F86303248D08F7594AE2FFF26F4240C1A6536564FC04325437627C804E5069C05759E2852D5AE2FFC2E7CAFE6ECAE64E22ADF663FD8962C9DA82C932F31539BF8AEE33EEFBB59B918F6C6E4099D1C7CDE7A4FEE3D4ECFA2747356189E16F838438C6523740E77D0034E82DE2E1C868D08E8B8DBEED96725C6D61C926F41E55ABD7873A6F242C00FF53F60DD63A57C0C65FD3E14267F87E5B04A1312E8945EAB4C37485C1B61879CD238380742A21DF99284EE65029A24801974B28BF02F6F0DDDD3B516BBCA4CA591B6C53FEC4B363CD634CCFC678FD4F5036EEFEBBF271395DEB4722272A1BA4B4F2D58F4EE2BE817E501CB262C918F91BEC9C02E6C8D4E697F282C34BFE68ED9B3EAF29E486F8850CF1AEA4531D70FB3C8FB8578F9FDC0ECF13D498B2DCFCCC7FDCAFFF124B58A60FC26069B0FB756B2B88EC8A4A90F5A2A625F82FB722674AFF9E798E86A2312C086919F6FA6CD1AEE32F16AB5144A1C1CB0CDBB1488A128BF058529BE1243FA63F0061AA41B894C7813C3CB458EE7DECE3071C8C5EF41895DAC9962B68284D9FFF798B95B57B1793B4CE5855E5A030DC9EB1888696CDD3C3A8DA23D9C7C16DFB0EF888DB99FEC08360A498C44D7098A2605345B33D2911B5ED4D507D5AC18D18EBC640A32793BB167BD0CDBD1AD091967AA4E45EA9F2B1CF982FDDD6A1C9EE55324C48EE03FA45EBF9597588C40DDD6BDB709D7F73E60F555475B460F7B0CBD3BC9D585C5B7BE9E6DE1E7C5776321211EA285F9FE1036A1DBA4AB9DB7B312C49B5851B38FF12EC1789F0F6DAE0F6CCC2DD073B4D0F73368231B0310E829907267136064A282693FB24A5E8D97006DB85470DCACAE09D0581095C03315C3C195EEFABABBD2DFFDDA71DDC9FE78DC70ED269959FE389D21BBBC75CC2F5D06FFEE5B00B4D08629286B8287AD514B390834D4359DE69CB868F8A7D5250A0812D533A5A4B3FCE184BEA06BBCB0D9B2086480E2DA250F4F6CD45288C5794B981D10BDA83D0DA9C9FBE1DDE83AAF8C75087EBA598C92A9F6251B69DF8A42C8709D899367AA10040E62B2E223070FA9B84B7A1ED84EF78A1C365346F25BD4266685AE8F23A4711B266245D085F8E3CDFBDCCF31B39EADE57AD137D85EF5DF0A719C2BAAFDFAF42F90B20673EB4181F175C7A0A080F1D3D0D1F7624EB7FE888342FFBBE83CB71143E708B057F9CBB9AF7EC68A46CC35C6E1A70D7A5F8CB1DBCED76D7AE3BCBA935C250C0A6892322D025BC43D8FEC3FA7821417D9DCA6B1CE2FE7E7767D61E73CD8DDD39C652D75CEC11AF0F8EECEE860C92ECE81C585E710A2CF91A960BAC49A98904C5A785F2D10D2E5D22393592A43E897AD0040F5971190441DD7216B789DFCF5AA72CADB2D1A5F0095A9BCFA8FC0A99675DC2F88DC24D753ED5AC686EC37D4E81CAE408A3DAA5C592CBF9567A446EFB244C5F84D9BC41AD3522E4EA900431507E197893921D40B266B86C06718F2A1CFDE5DEED3F1C2942B9317DC6E3492FD39D2EBB37BC6C4BE934451C3A5FA8236E6292CC8DAAE2798A221FC95150E464348EF45CC63F9092D5BFD809F33CB01E342A81E783F8499C02BDB87FA5C26EF13B7EA6954ADE493495294661357895AC57B081DAC9C1B958DD1C8F7E156EADF0247C60CD73F34A2CAD97C8F8D2034ABE10DBC5AB3B9EF11AC9FBCC8217862CF822AA24D077A652694A8924E2E836C9752E8B94B881D4E6C7C95A670CA6EAD88527BF92D7B875BAF45C3EB3AAE32C0B9E369C30BB3206B0C32C3491B93B14AEFBE0F14C7B8F68631FF1888BCD9BBFCD9F593095857F55F9AF30195183E3E8A9D589B15553CDA6ADC794AED429EB935918A8FFC8A86883479DDAB5EE70F0C1E7E30A98B1878160767C5E588B47C2947840B689480D91E364BAF30FF4B986A939AF9FF00B2D153C1878C42B8583258231C7092C016FBAED2DDDCD63CB3D517134112A033A74CE89F8E65BA6EC43F889D7F51716888D9F0D2F2CC290D34FBCF5C33F09674ADD5A702900357061DCA4E74B2E82D51D90A85F57C79CABF29366B057D2F248D9955206D4537919C4F48B8CC839CE377DB7D0AAB053D83C1A2A4331788D5A79DC18A75F9BFA69848EE267C71177DCB96686DD2660691998D49116E0867A0330A0E54B500C294DECF4C6B8A09875A9982C2372B24612284FF1157C4A75E1DB1168368D78A1D8E23292E86614274282AF92EAC9E3FE04F5F4AC6C890E4042DB4CDB6C9A2E86DA5D5B33674BE6CD39D64615156666797360C1F2D0FF0CA7344F693E42B1081D65E776FF3710F7F8BB691E46EECD4969332D58DD091EF8DE06E13BA2CBB0492B1DFEF1DF4946FC8D38096D5F8D4C5B97ED967B3E9998575448A7802628CA60DEA31F6D4BE9EC5ED06C9B50F5B5E171F0FA6AA19FB298A69106E4E92F4CB7801710F50CA7CC0796DD289A07A02DA6A0510DF79A3F76AC4C2F2D7E46CD15E7D5AF1449C65710B361D362D77C5ED6CDA8FC60C8D2435FAF93115329152916536EF3765FEDAA3FF196066BBE44CA6D45F02336C208F4C1A8C928B744B71FAB332829B979CAE32B5F7998E3A3519CF03C2ED1319DE79748077E82ED6F8336537537E2A4A137E6CC3079374BA287837D7E9E11123165E88A7FCDF68DC12C7F85D8DEF0197E97DADAD808FF569E3D9E1D30CA70D3EF37330F2B4A323E244F73CB3FBD18362D57309B877A7C78A4E0187FB4041D919442E83A4D58974BD8AA19FD9D4156F5AE58984D977475EF933EB11C2F16081C4CB266B00BA91E91730139D4B19AD6F2C18A45766627B97C420C6F81297F680BB169515852CF988B65561828336F573777D737FB37E464517B55E7784248B6CD12212ADFDCB134B83C46C1C98CF95FB75C6067A27438FAB0768E6DD4B34117D3862A5CCA21B6D21EBB4BDBDF97FE71C8D334DCB988F17AEE78921DBBC035143E248E1EEC745C03E6E1DD175B1AC2D8A42E205C17569148C3D3BDF2EAD2C769403CB56C93980F5FE2E25734190EED98E8E02339DE8F83D609F8373F9521B2DAE0E414F3EEA32E2373BF65ECF7E9A3CC418D71A9EF1C1A9F750BBA2420C1949FD132E66998ADB3FD94FE354E2035FD3C9A73F3D9ADB1100DC74D5647F680D78B7C0ADFDE96232EC1751F9FAD6255FEF05BD28CF429D315F6D4A34EC696F27A7195D981B48C9B8489A63403A02DCF54901169313AE06736D0DAA848ADCB431DB05F398DF64F16C1A65B4585DC1AE7213D3584A9862756E275FB9DD39620C47DEB248A578A932AADD26B3C98134733B4EB52968CEE57E03FACCB0F533E446BC8F72B87A614F493F273E196B0BBFDD81F2334C1273D27D8E851F85DD273D9D3EDCB886D298011651B0407CFC023B8785A2A6F42C010A7D6469DEEA1186067B3385533CBE6399598700D39BAF3F893A0A6CCF972482CAB4B0B1417200341B0017EE6F27FFAC51E067C15FAB8020CC5EB801E1BBA8653052AE6D730F1E3E49F423BF3A70DE96C595FEDA8EE2B0D0BC6B9456036FF1E041085E0D4FA15BF9ED27F548B75DD96F4EE911B357351EE2E16B8678B5848915CA65006A0CCD9394EB20003D976A0DE1DD81F532D76ADEF47943DFBB1D04726960E674188F3A5BF2441E49D41E7C8F5C91146C170EAAB94F074534664524790A60EA73D27BCE21124512AEA6CAFC674E2E27FEFE16D6E6DBB2D487AFC3B29DCC65BA50E0BB2810380B7DE1AF4F6E6B0F3F7F4F30B769B20D51D3077F723B6DF7CE52819DDC82B6EC053F22CE79A84E0D1B539B2960304F283818CD26875A561446D01B77A8EF12957614D3D9EAFDDDCC7B3EF70C0561DDB9A2A422B30CC381C974FE303FDF1308CD11A5ED5A5AB4D061B9967F75C026C3DE38076F3970994144CA966111F13C1C76AA9753CE588490520619F31B86882670076600633855ED38A9B14AA792F4AC0C15160D547F267DC8EA8B44617CE6E0F16ACA3BB58E22C2D024D3EF8A613593F50CAC95A501B00DA8223745AD11F9C74F7A85BC7AA8AB621036AE644022EF7DBA6C2FCCF08E487C64928B8DDF54D3AF8157B164631A3A0830D26C20DFD0AFEF5AF30EBADD2A864EA3F99F32BC2D99F849726AD445C68718088AFDF0DA43910CB406627E425DA136066CDE45CB32E2AD19992AB64A70334A5A78C31A08E2DCD3233BE097F81060471C30D985CAA01905B1D0CDCBF203BB0AC94E679CA5218961D979EC0D3A2A8F1E917F2C42483E42E42C92FCB2E4D580A0D6B23959197F24166355FD240CD372F3DE20FCCF3532329AA2D2772B66C183D0019A3FD77BBAEFA1645E4E0C3D68B8314280778ED4CDC6EDE526D98B960C10524967B42A42B229351AC026400A986D2D48E35F7512FE9FBFFD26534FD2852F1CD2D46D046DE732A2C264F5AF7BDE15EEF3A59EAA2A5F220FBA7E81023FCF4C4B73D6E79F7784669B51BC5F88F8D3B66A5B2F26B98ED96460FF80F3CB4095F7A38EE0D9ECF47CFE56DF2944B4B7874F01F1B4EB67A3B35975C32FFE0DFB7FB96BCBEB845AF66E74059DC88FAAC4582949DE01022A79AE32DDBA77AA95811F554CB5556EA8FCFB93DD4E8A04185E2BA06F950233D0BDF5C08B328C394D677C596664C5D403BDA45604AC777DB8AB34E1AF1D459A5536C49D314774711695AE298D2A843AC838F0D9F34B103C32B3CDC9512415FB58C2EFAE0D35C7DD2CABDC0394173498DF85ABEB11D318BB09459081092E567B516EE0322EDF499EAAC992B0C50C2CBA8EE2FFC42CACE5CDD250C2A817C88EE2399554FF347BF5BFF8FB51C7CEC8DD6E97AE3D2CC04F4D2D3A0A5D57A2129BDC5B50CA2985E2D6DA03B6CB286937FC0D34E5BDB82DBC668B346DC8007D7BD065F91307FAF3B434312C117F357388C6B5750F36DA439B3D3D4D6E5793FAD17F4EAFD9D62DB3F6B4EDC985D4C39FD8F34ED460097C1BBE329F061ED674CEF54AABDAD5DBD95726C77AC6F24EE67ED41BD496EC2C24A23D6B0EDB1B5D7C6B44B4B56E07359DD6B052E3C8C75DBA1CB0EB07116C21B2C3DC03EF60F769B61B8C40B84444E571D0537B4AC4631424FC2AC1EB207DC47773BEF2267A11DFA86DD392EF783711861B81AFE42DA9E69FA6DFE84A6640271E40CE44AEB99BEEE2DFB4C759EF63967094B938832DE2509A9B1629FB7DE1ECE41166F5783FB62E7771E806238BC44F510341EBAF71AB3190DB0631566F33DB97A7971075AFCA63CD7E9FD6C47648BBB236455F11E5F18A86C00FDFB2A4B1093F5DF213309A64DAA398684D9BDFE1C4B76109980230465FEB97D481D8753972241CCD2EF35AF41F3BC943D2288550419698E21966BCA5948ED4820221D7C30D0B3C01D030A2A73503D34D1623372A4A8D8EED08F32BE985A979337A58693E0634513642BA7E1C52FD0E4B7DAAB83B7C54C985DBBF3981DAD1FC54F7F62AFB12A30CF4BC44300DC453E5B3D710A350582BB8963476CB0C820219C2BF07C2DF4C8F27A0C4AD65E2CBEE56A3323E90EA9CD71CF00C1A39E3A4ADDE0D9E9E59887A751C9BB65AD7337B86694C311C2FB75FF567961DE80E213C7F6A36BF6DAA7D5EE471A520D717F05FCD766EBE0D48ECDCB765C888745E73B84811EFC5D9BAA0316CD9E315CD386B251723BC4064F4FED4DD7F70F4A58965F059E63E0DF13C1B2D3AD06D0B32BEC46FB5E6EFCAA10A9B2DA293D3C7EE848636368966D9CA61B57B9E9F41FF0C4BBE9F8DD9BB991B9D96CD32C2D93F3C4E63323D4C51D9DB8E0455A4AD317D816B09F8592371D85BA24EB49A90835913245BB7003955D6D5D6B6796CE3221468586D06E26B4FAB17D09C525F8F2AF25371C8A932F228455829998D590A628CE314AD8C7E1F7E74BF4EC7623ACFE749748A22BC392410B38812E7C58A5E98559DE10AE1BA66F457DE2425B4FA579987168EC79D6D235CD78D26378C18900815867282811D3A5DD7E3796CEC64B4D8757012D63FECA0099A57F4B1867D0783A9ED9891C9E9212927EC6DD46C57EBEF136526A4800B62A4A854C46573B51E5C8042B9D9F3409585B52660D3B5E49302E581C88CE17B5187273B2621D75F246E4E08896D4204DD92AA7E9C2673BDB90819FDA124ADEB7DE9368DD150728642ECFA24856514ABDE4BA5DDB555D96445CED7931139F01E060C56EC48868443D51D06A21B5DC031871C3E3305A3C46D3059EE862B6DA0432B7D81F2DFEC9B397285B0B32F24B6CFEE219AA95DBD18F9B93A99FAADD5F505A1FE61ABC70114B29CFA8FD9519543E6A4397C8240D1DEC0CB5FE5CA8F2A4A256B5CFCC7DEEE10AACE1B0267C59745DBE6B16D133A9391218B3170CDC408810B24AFD5DA7A2647D1798B16F776D9AA2C95B53A6171FB744DF52248CD3416ECA68BE0B403EAEC235D87F9A9BB586DFC1906D86313314B54D011FD847E81C62B972D24F0AAFB401F6BFD328A7E5324057EA94D4359234DDD28CC944BCF4A3EF9B81BFB396F6EB4F5BEC38913CFB07AC208B65A0FCD889BD0928D1F0A40241375FF5554150B5647AB536E3C71846D43E194A7373E28F04A5F95E9ACA2B6E2D2270D7528834FDDB7F71E67824356E2B46DEB6272EF93340E6011656C14115B61C9AC7CAB0739129272E426BDABEA73102F196A562F7DE7FC18D4B1129A966FB80761E400051A45B991A144E5ACA472414EDFCBD1FD5766B11A5451FB98C475D98757337A98CD7AC5C90EFF48C3082F79CD80F103B5F419B3490A80AD02144E514BF26A43CA91434928C1206E6B51F374ABAACF5A5FD3DDC6C00B8A79B8E2EE7002EE312A33742135BC32C8BDEA8BF7BA7A1E01FC2FE19732C40C6A87845F71DC6C814921C35B40BCE30291BC404EE3B10A01499BF998A45DF39D941450A80106C48B9ED73B7FC26025C6E0F241D1126B5455ECD119549F10AF83C37D89648BFBCAAC1A655CF5F5A427B698644E9DD1E44E6BA8EEBEBA4A9396F4CB045C5E7BB10C338BDED0B71CE0AF787BE723F95861F9F29107EFFFFFE429592449F94A9FDA0C9EB08D0F3AD0C0C66DA3EEC16D167768E33D044D85E4FACDF45D424042707CAAEE613CE674C2D3ED409C4912A049D4B478BFDCA02E97208BFAFADB0135CC3F6D707E07FCDAE452AC2801F2B851A9C23CCDF963A7728D31D523B585D8823D7E4155F8BDDBB017AE7D298BEC48D60C0A51B9D9D01E5204610032151F0C0827A4128BD6620647CA5C5218FA2E0D8731760B8B43673EF2B35DAD0E0B8D75B9DF412CA087CC1681B0E438733A08AA47E8B5DEBBED01757BDF3B0E84B683C89710EB18AB554B155E7C2B7BEB1A0BEB20BE1EDD6ECCC3BBEA5183EE64EE3484BCD9D499FC262C7884DBC1BB381B5170993686C4FA89EC41A5DEAE6F2998DB5E0179A957A0D265147777DDAC518CC4C822D8EC39FECA0BBC0D2585048CE0C0A8F98F28C37E891EEC632EDFD9C19BA0BC20DF434180C912B98D0D13631926DA4BB087E47BA663D0E633A76BC3A28FDA39BEB4EF1F2198DB269E550642D413613269CA9C40D2BF4A20BC1CE4F6D2BEC2450DB8727E498E6565A2EF9BD9EEB7FA48382F665C528EFADB3261F84E2CFBC8C5836E4D5C8186E29615F807B83287F561ABD3F276786D40AEBEBD971C6F90D0F9FE46EC637ADCD9C479EEE958F8E6B1A7996C434298B6D5667F07C238684455F70B647E628B6CC77A57685EE5B3F7BC1BB14268A80351125CF59D189E3C19DC28D63EAC212782D35C57A4E825B4B93CC8782494600B60CBE95CA8D107EC45275B088DABD7186A951A4F0ADD57854BBA4E5A04F11814B25557F53B2EEE6EB36C1522155CDCFC986C5B5DF4F6E96BD751D898961310AF7986B063A6F39DD1D2DFD240D85CA565BB29E0A15A4556FD087C41DDBC4B6B970150A41AEB6970B48C39749CA20FD29DBBA23EC3FCAE7E4B8FEAA06DB5277B98B713C53D16E51C707F7002353CB166F605B229977A2D0F15B454FC338CBF1079C392E4ECCE83ECA17698FE7C4D04C4E978275721C269E9955498EF9CCFBB853B3AD3AAA664EF05EF2B771E950C23F7C8A094C2F394B390795BAA0A8869E9C086B24D3D7D9CE8BBF978AE57FB80A9B3481A4C79A0F32DD9E21B5F24385067B3A3AD4473E16784AB8B6B9B43E95DF33FB3B25AB0CC79B215DF200A045195F27367E880ECE9215E9BD1FA85A2D87C893C4C49A7D07A19ADDE815A0435AD69697BFD49A77B8CB77D462AA5DA93D12CBDFC2D79F4780427B0C97B90CF3BE2A581CC15525A8B486D432866B347FB1E0F91E1514703119E54248CF5456DC5E6B8CF8ACCEB99D5198E4C8C07177F4345E8B5FE1E2028CF42C334CE945CFBA0BA3A8E78E1A08A4B3208E33B8BC8F3D06DFAC803794992C71618AEA070ED4BCAF155648C72938B2F353EA68CCE607A5B2D6952352D973806812B5877D8DF35D9CBB79870CA745E5C27136E52CE29EAFC21547D332FEC2D46F70F6F98359B33DEAA312B61B995C015940FCD16427ABED3DDA8E4662AF119739DA7627DE1F38DF6C1F9478CF381A463654516A0E6DD641277AC2A0B235173E6CD5487EDCFD2D7B89BFBA7AED977D6152A184D10531533076D71545202F49C5F381CDD6A80FAEC4CFF19235BCF4AD9638BD613180A96D3DF7F9B3AB5E9C10EB6F9A4B3A7205A0A51D5377EA8C9AC8F18DA875360FF2D67BC0A630B348A782E20FBB63C7061695F9B505690FEF5575D66DD65ED4ABE30AB8967311D8FE9A67B13A62533D3BC340ED1A50638748DA6AD63C1AE2071BE84BE4477594B3D34DC24A43F8FD01E08B2E76D9BE4E72069FE8796EB15F1442EF686FBFA588CF79142EAAABDF4DA8D26761D97066FBA719DD83C221078A8FCB6FA8532633FEA9DDAD1BC3D71E3FD3DBF351F09E3577EAE8E55A48841C23D53DB3BDC3A7C3D4DF635487999E8A3F5474CB26C5E1325E4D32B0D0408269CD687E9BFEFAA28886BD8A02AAA6ECDCD2240505E70E30473DDB811C7FE6F207FA381BD028A0D0522B001B585E61788F68B9982B91B806728C0BEFAA443C7EF88A4858F3C61D8184A9A1BFA96EC545C0DF3C4562D9C28D7C16FF223D8381C93FDB48A64969512866A68810036005FD2CEA7B733D5B68DDD76ABDE5711155A88E78542E36FB4A1C2B809D8A91826281B0538C6BE1EC70294C09AC40FA5CDA7DB51D137B9A6DEB997A9CFA3FEFBB441F72BB45FD07624EAB8833D8B55ACAF8B0D07EEC2C2E0A74FB71144DF44778DF1C218ED5A77C4AD32152D4BF8763F8DF278FBDBB31493D3015305303C63BA5ABB08DB29BC17791AD581FC03AAF4770CDBFA3E2A4E3650830593C10DE54FF57735C519FAE8F3C80CCF23B373A70F56648E589BD1121DE0AB5AA53473F58FDC036FA00228E989CDAC1868FB47535E8647B0EFCDD096DDE65F70E52419B021B46AA1C58D18BF6CB373E61805E5ECF2F39227478E3EE82717D60986A2EAE901EDC0CA97DCDAC80A9ED943B2F591A81C685308744A7302FB36AB0B4A8FF87878050F6998740E2262AF2D88A7BC8EB982106F872DAC50E375CC7B0C084885965D97CFC2B376A565D90087038169406E98E131DF265833792929CC4F90EFE7FE8950420528531559634E7143AEF3E3616944AA06B86FD39DCABB81FA2439A9162EE0E91DAC971219E2C73F5AC6DA07CF7558BDE3AABABADAE9527BB473E981C950739F85209AD36BEF32F0C9E5007FD047147D6298741CFA223CCF017494998B38413813F9DBB5AF5469D1C5027F59D24699AC4E498B4F38FCC4C1C38E5D0153E89AD1F51B87F97A3B921DD02D90AD0750B24DC8342F3B090DABF06875A64158D4775A8C3D8CF0358F160F16B3A4CF0A5DC646C00D8047BB1F9638F03D5A1A84A28928FCD52E0CB00145B8F5CE6A821ECDAF308CE5CFA1C41BFD0071DC3BF7B2111C0B4414888911CB63CEA64D064487A9DFAC401EC2CC01B9F709BA5244CB767CB27CA69E1D3A64FC586DC56EABA7777DCB12CAE2E2E30E7662998FB8B449B0EF6EF244E1AEE8C7A1EBF685F0684E9317E579906DD56B8A7D461CC69367F6CD017A26EFD2ABDBD3D99A3E8A85F8C98E3B1F9F362143DE109AE847B31285CBD6B9A3A4F46708DC262EF8C6115C134E8C5BE9248523659518360B198C7618BA059C0A8F0740CAD4E15AFC84DF7E016AFBEF983BAE8F87B0FB52EB0F946EA08671AE115055C3FFE07C569DB6DA43445E9F563231FD1528A492F65D6C0800575EFDDCF4AD689FC34D13ECE02F46ECDD24BF4D5ECB13BDBEF341C8305A86E4DD98E33FAAB27B037A970F775FBBE0DBC23CC590C76A8D132605ED1185981BD9746C2CD990B31DDD6381ADD69DACD2136401E7C197A94672A5D042884F68FCAB5458D48F2EEAA56410EADD3D172E57DC89871B5EE88A410CA5D7ADF252002B487C5BC8EF3CD03144C250E6432638558871BC61D5E348E25AF43617AF5D4A3E6563E8499BA7AFD1835869FA496035000867299C979D12D768BED5DF76C19A594B1D90B5D2FEB3EDAA255965BD78DD72C908B68B1D8EC45AA6632CF1C95F835A61D86FCE02AE40FAFBACFEA7D929824AEFDE34704A50ACCC39C3B168A6798A4272C6FD3E165F9F40E60E12BF88420EE3471253DC714D2D12F9120CFEC23A73C2F4B087537B8F6359ADD70835F4F741BEC4B0BAC1A617FBEA82A1C856BD8EFB34F93F84678B43618471E3BFE01DF2331212B8D66CE126C5E02436A2E84B1EF792390146BB1E3A20F9732F87431834B8D80286BA809521E447DB607F26341EFDEDFEB3A46E6F20F338397030F4EC15B3113566F4871E195488D937E4F2AD3DC75BE6C8FD2DAC9E3C171D474BABD7516857DAB383A8DB41B6D952AD01FC9CA566D0110EEC46001F3D2B40B024EE09D86D870EAA383FB78EDEF8780BE35E183952E1FD10372868DCA330F4AD458C769579A613A2367D4F06214C4239D0B9C1321B1479917E04EA4EA65D4235298F960EE3E0CEA3818EEFE1B5D94387EE2A8B02669119966E2BFB0FCE36BFE73061EA9BBF09298B02185CF1C5ECA2D5419573B1F7FE8D3FE3E1A1BC44EAC4B602B766720E717D657F0BC29014E9E5C43075E74DE0767D6578A8DAEF80A4A10E08895433CE5B198F895C1F406D9F1428C0758B888493E16822F253A32F39D1F3AF4B5697773D8FF9B43A2A88DF848F45703C58AA1E61FB8487CDFAD137E7C8F45791E9B87117A256484EDA1AD4DAD01F610935DD4AA1C17173220343FFD70E53D474F4D511FEA5B97F302DAE54465C5A481AC7CD96890B27D6405FB2BA8157AE5F842D073A8155C2A843062D5B6673FF82B6AE5349C0AAE2E429478A68FC8F528FE3413F5901B3C331CE34AD7EF9E2E85AD9EED402978FDACB2D53D4F7B01C85F4D6158204CABDC4A3A6FDB1E7CEF7E6E05A58A5CDC172FCAC695D605CECFC60F952A934EE3896ADBD43DB96131415B0ABAA812CA3D849A5CC11171252EBBE320BA689CD453964D5420C42A6ADCF6C7A133E35C96DA1FDE67B89A0D5F967BC3EB09779EE1AE78AB2051810D5133949C1634E62CBD33E910501610E8C710A55D88E35FE2C7CE80CA31614872C9F1D409A74B2535EA255DBBFF5F45F7225F246CC296BD580D4AB5FC4FE8B78B1F62356A4DDCF6789966605F180DBBD2233E8A75C277D9BB267EACF7493C8D0E61A51DB30FDBFD495182CEE17F6D4270014379EBAFBD343EC6C5AF9862E7E500F6B37BD000E5B61E5659F5CF7A629A248A1E8564F17334F90B686179051E937088FC1F20F1D5AD15B8187E9AA8F11498261FCD50C328B0A740A2A73DDA772219ADC8AA6F94BCA70C06F0E457F19A4054F3F96012256EFBADEDA186F76438C088D2AE8E975CCCC0CDD31482234026CF860165A13522C3077AAB904420FAFC5D2159BE05E0217C3DE557AA44DC11B412938FFC53CDF4D83ABDF261B8B1393A017EB88F449F4B0545C0706F17C2E265BE6EBD8A7FC02C044B6D9B3B068F554044173F0BBDB1ACF82D770567AE7EEE432427BD14875DDC9821C0ECFFB07EA472BC00D2FDFADBA1567307060B8B6A287BA8BD72B232C7CA7CAC9A9DF6953099644B9824EBE6686CACF32A4D520416FE2B07482E1216EBA303607F83B6974DCF461D0E9D3901437FC58BAFAB2C668755751C5C5C8F632DC41FB4F75A7A9B8325863B08DE4CE6F65DAA80ED2C353A62E654467FF7164345EE3A3D6480A14DAB149D76520ECECF6EA976553722246523B9A92EA38C97276CC48B66E15960F2FC748681AD1D5BB80CC0ECAC31EA1D6B6C5CFAE0D56CD8AB352FC6D48143FDD48049DEC8D9F07DB0A8EF59D1B06C08E78C29FA660C6D681B7087CEF90F318E814C6DBDCE053743339B9FCB62B2289557BDB8F139720009862AE6A084C70A101A506384F5EDF12E7075D368BCC4F5099C4954535C7BD6CBD890E5E2E0FB8B27C98EA36D47614F6337EAD2649E965B0C5ABC8F479F3D0437E10514D892936E4BB05852ABBA8A0A125774C60C8D70AA3B74562BA600F70C1B97F1C1290D15DBF57D99346185614FC265AB754B43D580F6CF6A78152047E9EC2F93D5140FFE50B0BB1F9794B5A16EE7AB7305FF969FEB5D1A93F43E704B44635FDB73D31050E0CBC8CA9FF3C41F7F36196AE1FEBB18C2A5F72BDFE69260A0517D86C522A005FE2379410283CB558D0CFA424764BA10A2508ECDA941B23DCFC50B4B4E1D13E9FBBFC70F9A89E7CCE29B21CA1907577022C695DB72C38AD3FBAF9F00D84FF0CE5EFF1CAB97500F833DF1D29FC08C06C9B29689D7D2A50D8878612D1E805B398D40CB1D80782817DE18A7F936D9EF8D83A481079B55E5BC10F13887B8132FF6AD461F666E91EB64262961E05C979847250969740ED9A7166E63611247ADA568424E5BAF6CE77AC7463CCC9A8E9B826B896223796B41D84DF60516FE5FF7F85623D7082A786B7ED8DBF1836E4999E81BFB237B22290F91CADCBB2C08C9733ED018563D64B548606CBE384A48D020CB805D3693BD6651DA5336A15A71C16597C9187CE3E530700A7780F54814527A3CB41B28FEC68CE5D24E5A5840C46FAAFA96F86B5AEEA7EDA8501E1FA3FB22BC890D44A4B1AA24F2486C90196396534F68C9C48D3C471BB5BC61292EE9D936EE839471C26CB603F3D53AEA83BFD07C12B685255D6A028CD4D4088B8A69C0ED4C86128F4A39735855B04C0EE000A521F1A754D44362EC5FA5CFB22F80D75722736F27AD0F7CA81E532C017A28AB7C083F98238B9D7CCB92F46DF888D839900042C72FDB707DECA62F51DB3ECE470FA2CB58BBD9E93C09DB6607D0D47322836C811F77468201462EAA19488784EA59DE6AE897BBE1CE4375937F101DB75B050237EB1DD711721DCD05EC8106579D48F7390DB18BD14908FB50A7823713ED0EFE48E2353A9125C45B002D1A904BD00630851D4F0CB5F1118D3D3533A9D6EA07D0F14E29DE51555BCE997E96193243B47CECA5E1A1460DC3490F06308C928E4B39372547E09FE2A64C03EA7571043A8911DDB1D6D2C2B2056FFF52F520F05A16C36E978A4D7B7A6F0E1F0E67727C328A53D3F28969B543AD0C6282407FBD81A57F72D9730D63A69F51C1E777229187868E438193E8DB00C5B67A63C478D0F5970775FC4856425C3F3A38ADD59236E9AC33DCDC8F49CDB4BC1E88DF33D032260BEADFB6BD0D567794800191E3295408F8CC5CEFE680672D633B03DFC364C254D435F0C666EAC16F339D9B51290BE646AF0AD172294ABB9097ADDE75969751E2E5B09E7F9B3A8862B3BD454BC7B5C42AA0CF53CC1A9C32F700CC264D4F395F45869AAF4F25DB36FEDB8C19B8D3489CF7C1FA2F924A43A98ADE55B2D299FC0DDAC799DD62ED6A10C954A266E0B80FB589138BFA98CEF25C9A763227D2716662623E89A85A1E92CC3C127087473EC2A64E6A72436DB44C468A67834EF1EC876354B525D46ACFA8A9846FD0C50A4064BEDCAABC06CAE5F03BF76DC1213AE4CE6BDEBAB29A457EFDCE9424C433D507EACFD1A19E73C04FEAFE7B96554B7229D2499621D0F4B255C34A1D41B1DAB44F89811D96EC3FC31CBBBC4E35FF82FBFFE84A2FED78C870111EBFBE71D0F14F12112A088DB8540B5578B7D2F478238BC1808D0A3DCE1DCD5C4BC767A4977F69FEE36055ADACB9D7D689B95AC4FF2C325D4F708EBC96D0CEA3BA1BCFBDAD00AAC13F92DD92D351D518961AFEDC55B2AC6D6E28DAC39C3C5DE994DE26A767E64B460D08D87439ADE5E901F1F16467104CEB73DFD13D78080FD9F1320E27A26EFD15700CD8A2C6F19BFD965FB82CFEA7002C0FB54D6647F19103BFDE255CEFF266CB0B76DF52DCB89945CBB9AA0A6DB37AB48885728F8DEE9E153208FEF6A871A185CEDC813399CE83FAC7D7A0DE17A6AF789392E75480071A5FD03BC0F9E395C82F72D433349F08BEA5831D3566F5A46D330FDAB265CD739ECEE9D460DCD5BDCD1D10E6567AE85B9EDB1880015C7698AAE6BFEF8A0B31AB5A98B14F652C0C8AA0F2B0141D386998CACD8BFC3728C641F865AB75F1EE80E0E0F4B216CA2723953F8A6B1E95E86CA513396A66C6D91D12393A997ADD7FF4149B3640DB7F4CCC927CEF3D9D909BDA8E2396D90EFA7699FD3DD233510B394ADAC7BC7F6218F7716D9DB6E91C4B3D38DFA342E46B310CA3B26761C13D5F2E99020AD1A8131B44C7AC1B48FD8EE242FA02957038201C45DEA795410A87EE97448171602B1A629C43767784E340436C14D2E295831EDD2EA82A929963F39436A2125E866E98E26DCB4F6F6D9DDBED5F2B13B62001A52E4AD49C0567799A5F4D11F3DDA976431A52B38837F15BC01E5E4F113CD27D50DB3BC1ACD2A42E35AF69DA7852D83D06B4E13BF98900879491A30D8E783D32E5252439D6EC0973FEF6FDEE1DC6EBE565A5EF05C2513A7B290D52C9035FC5BB7EBF5CCFEEB5D483EF583955D5939DB34FA5BBED0B7627C604A05ACBD2655883C6E686E7BE74B4AF5682834F9888056FD652462989E1B9B832DBB291D3155A65B5C3352329197ABE37E4670A2ED90B5C5FE2E5AE5FEEF0E1383B397536255124A5A676B8CB75A5857F1277D93AD9808E996419D40E1F0551F4DEF63F605722E1B0CC907A322CE927F8CC1CEE496886D50D35FA22544A95F07D8C33796917DC2C2478474AB6AB956307A8F757194B698C0B89D592177D8EB35D4F994BB8D555B37C7E13B50FAC14C50B65140ABFCCFE1FF44E257D9FC9B84240E98B2BBD875123C5BAD02289128B8BDEB1805410BB90A3F727A9FD53D849F9BC3B624CCF1D6E0E6A55F05E5C08E2A5777CDBD5472DBD3EE89099F7A00A9F35EA51CBE01FFE600B5C9CC8B2880309D88F028A88A8848FBEE94076FA186F5BDFCB5F4D09948113E27D754BD1BEBB06713E0FBA44AB3F92DF60345833A8506DF162046CA4E32E40AC85E370C60E505CD387680C9DC765386FCFF66869F8E00FD51A65432B40CCA2173DCD8EC23FF1FA8AA8D5EA8BEEBDE25E92FEF40D3CB585C84428C766185BE2132EF86F97C19D10611A5829B4A03819CC64C575F0AF91AB6E8A7CB8DC4753A3971CA84D10CAC122AD260FC2D99947A444A97055AE57FD77B23D21BD0852DC08290A679A3EBFF5AF341C29E411E19362E49CE49D98DEDEFF7A475506DEF6160C76A3BA5453911DBD4598090FEDA22056359FE472F2D9F882DDA0CB328BD402C73D63EFF115C58A50BEFCA062B1A750BB64242D7ED934A473F52E6BC4D6CF687CC6479556A33E239C4CCEA244843AFCBF9E1BEA6C977411A142166A8B5C2BD4ABA76EE8C467CC6483CC5FC183350B97891CA90749CF0F0371E34AF156F11056A1A521054EB7CC0410C5313C3D61132E59C78ACCA416B01E2A381E663F047D64244ADD142FE358263F998AD81FE9309622E1F8D0E46195F697631857B365E3559D5552AC4891FDA31D8F950F9B546B4C693C915574B0E06C55FDBECEFDAD99CDD025FB3F163256C68C49CFACA862AF66CA81D1AB420B497F83D265448DE2050741A814DA0C73B9FFA46D2121177F938BE42BE2C96D5F2C586FE33E2AD2B589B27644855F6053BF1ACA18E6BC8E8625B42BF9A1C72298E68091BAD3A8F532E6E5612F55BE38D07AAD0F34BB606C40474859D92BA3BA53F1E9958795206125AD2E9A069EC182AF31EAD0B7512EB2DCA01805B5175AE4FD3A932ABFC002C571E6641E5DB4AA257DEE482B3871FEA68057757A1AD8D923B250B8D89391E9C66495BAC5AB52211AA8D119D0AC55EC3E94676F116E4648CD62E2566D17533BD9B832DF9F03A65517B0038C219B82DC07A4F100CF202A10E84D7FDA6607BC41E851C2F5D29C2DD0F16AD42E7F0D90106EC9C9C62C92958CADBB04CC2D19D884B363D20A1497974E8684F4407EBCC15BC71EF78D6D216B3B451B2A3D724429CE216CBCD76A8794B24EF2C3D758BC4F3270C9C5653D9AD9D77CA271B7F546FA4AD05BB72D9BB65C50A3C267E1F5917385C937ECAE7222FA2A371289B4688232C5529265B813E921B569C96279881249AC1565362B575CED533AFB30C03E3AED87F96C0E3CCEFE0BA666D91384F17C430247BB4ACAF5DB9C39ED41EFFC065AE8C4437D7CFFA190B5C7892BF7DA5032FB29334AD01F164EACB8E001A749D63B5AD27CA3A4020492095299F372CE1F3402DF3057FB72BA75B5303338AE907DB9DB31056F598E3A32537807536E68DAD12BE8DFBA49B442BB4C3DAA66FDB1CD66D98FA5F29ECD67D6FBB41C81F5AD9508CC6C290C91E009AAEF44C8756E8BAED964F224FE1F6D2BD02B330E418192E716D036E4F7B8EFE932C442C4F6CDA26D794C8A6B911480EF5D2655CCA487089470C48DD3FDDC0F027F714DA4E14017AB5144EE75E7C87435B315D61D7236FA0EBB81B4207B11F43D6DFDB3FEA6FE8E9717F002B4C0552EFD8289758DC92679BF28FAA032019ECF14724664EEF6D6A29D39E9B380A9BB3D0FDAFEBCD43213E47D98D7373A532AA0BD44FABCC4D5A3BF4CB02E1501F4CE69E05153B0F22BA09BA3D37F92CF33A0307A24DFFE1A2430CB798897B9D77F8608ED85F71F172A72EF3866760C8ADB5E0B77CCD58A8494C48770CD657888DF216C1F393DACE0C68DD9DD621E52D221F3E89601FA9CFAB04E533AB46C533803229F80EA987037D97ADE9340F5CC84BCFF37F93DD1142C19B2A1059103AFE642737966B05266222A1542BFB699D3AC69AFAA4EE1E1BFFD1B8521C59197ED17DE1F1B88697ADAAA7352DA3564820BA8CA1E40B64FACBC1C5564E25E01435A535A7F1A8FDBC57E85F374BEB10E576E022D79D67F830D850C11C682D2C962F0B3C083DDB3D4C95F26B83ECE438ECBB0B0C89F94039AD21B65379ABD0181B8DC88961AC9990060A256A7EE7CDA27C5F4A718524F2EAA6742F7DF37080CB5CB665875D8E084EC8424A1AE0C0B96DBBB844B3DFED6AC0BD8FE2EA00B91E919D4B7A600E27C3948A4ADE23703C61D01CEBE04DB7ADF50EA54DF5BA26D25C99AF2C9A9637630E95487F59BC40E6503F1B570F0485E6BE7A0A662D3D83EFCDAB1AAF695D3010F810CAAADE589F6F76BA5B4EE43ED39B39A19CBE7040CA7B52663D146A4A37B8F3599979E209AB9E99E0760F24711A7F5C6EA4778EE8EA0691241D7C062B9F2C1E8F47F68613CB2402507296127C996F01AD7035BE4A7B013E2F91CBAB0BA98C97DA648A2D086BFAC033D93FC983DC75B28D7E652FF4B138FF52A877F00169ADC706B55F84674DA6A369A14042CCB42CF7F1D3F5986981A67666FCD69ABE367CC2BF0DDCB9F044DAC9C2EC95FAD266D18CC72E3F46C3A08AE22A5096FE7DB9FBF202AF06F3CAB1336EB9EC9F30A40887598B89B49D0899AE4DE020E3735E562BF34EBE4F6089592C71E84C19998A155EC26396F1C5F0DCFD646F2BCAB5781E83CB773F0081E864FDA6D1AB1349FF9078C5288F29E6518C52E38341211682394673CF497D7819B11C9737564DCFBDFF5A32EB3E25A96EBB0DC4943F4BA890A86F67522FB7CD76913432418B948A4786B6C4CD69168E6756BE151FF5338297B9A642BC5409BF054368ECF21C6C7BDEB8307A4AF4A33EAE170A254391C2368F03DCC64AEF914D4332650BEC614E99477F86BD75FAAF9933CFBD485C38B9929BDCFA668806856549B85ADF1A629F799D911CF7F03FEBCBD6E0F7B93DB1ACB0454EAF6194FD37C0B6C81806338A062F76DFA3C8E2FF6AF5AF6EC74912F5BBD0F7E53FA5557F65778678A273743ED6A60ED635351F2E7EBEB015AE1582DBAE15594BCEADCA0250F8D0EBF32209D626C113ABD6D5A76A6A63944E62C2B59671853781ADFEDA588744CE0C17846BA75A863AE08719A5E6AFEEA394E105DF7C73E16CDE8BE89E6E6F46CD2487537F6A442E180E7458B593E74294A385958CCC10BC2F435A3F8085DB47713AD5167BE8166B41F8A781AE2E9E706197769D3AAE1600D892BCDB8A0A52E8397159EDC4D33C4533C76814CB4DD247C949D1A99FF2774721CB98A832C179ED10EC5A0CF29DA7EE720C338FAB580E1135E071E261BC5863B089115828089F25014C106FA55C7EA29C5A1AC96D4D751F61C1E2D62A065E82A678F1517B14B9A49E076CBF5413AEBA50104F0CF8E1C38A03740F8E13CC57BAE640F8A022DD66EDB9C2AD6CF9855D818413EFC9533158DDB7B981F3A3FE6F0CFB75D495B6F2ACE41C0F1B65F83B83A71A772B8D3DAEEA44C18805BA9417D30104F3716F475B7D662981209D856B6539C4D0C9BD472A4ABC8348767FB217386670BC5CE1198D5E0BF5B365830AB0EEBBF78F9CE2EEB1A8D3263ECA5983EEB096C270DF7222A4C191EC1730800D48BBEA88D52F5B0681F55AEA50368BC2AE1C23DF021A55A54BB0427DB078789878CF5601BB3CAA1D22141DA87FBC953874AB1579896D396E75DEE2F1DE932EA206A15077EF41D3DBE950B6BB28B3D89FCCE48CE42D073E31397AA7308046EC5B2592410AF7807B11F1B92B66A1E615C7ACE0B075469B3418F85AD620AF827BC289F957789AD2137D09B91050C4C8622A17B7885BE93E449A3DD7AEE341EC61F07BFCF04E9066288CD7C074EB9C3042B7E670680D26F5F529A7B5E7CB05B1A1458ECA49F402F36BCDAF3305DEE845CAC734E3BC578B2B19FE655849CBC11845C988D6DF26BF9C2D600272E32B2001F33D87665ABA16EA670210E9D45FB7A40E060DA8B0D76DB97DB2355EDC721944D4D050626D85F917A3ED151FCDF6C52AC54AFB9D0B5F6950951F97400CBAF239B8E77386737D10849F80C704404F7960510C71FEF9197C38E9F7482645C17283A86ECB3B42488936C2E7F50875FAC1E699B10ABDB0C5571F1945DF48FD01D391937A410422E1F2E3117A42940CC1E5E3F0EAEC8AC54F78A07649005379A2CFF0CDE1A6B0B922616CB19573B66387A6171DD3CD6BCF7FB55E8948E2373485C8EBCEE47A100AA09B9D9DB468E38E5828601BE05F623E1C4BBB5B2F9EF7B464E5A057BD57838508DEE1DECB2A3FB6394F6231791BA57BAC54D162B1F0A41AC3FA0361B413343F0A901BD1116A66F24F1560B81F13AD35F6AEB8991FE0DDE0B77E33609A9960FC52FD8DC09AD708E850CE8A52FDB89650B5FE4C56CA676B99BC604D7AF68205BD2076472085A44D9E01AAEBED160E6B594C8208F0D2A6F753B9AC54AB5E0DC2D6C8978D8A15438FA95DBFD481C70EA1ADBBB2059CAC89FBFABBBF021E27C8826D8F3ECFE67148D42B619E7C13FF03388DF548991902F197571E62ABD14BEB1F5A158FEFA9264EEDF3A6F5D1274C3450B65676E2BC93708916BA32F8C0D884DBD037E94865CA4024AB737762A3C156495847FB96C6CEF46B10B16560E3002C37753B3F1CD5F4355ED32BF5E2188660'
			},
			SiggenCaseItem{
				tcid:      28
				deferred:  false
				sk:        '4413FFA029DD213883F0577CB051D5DA0BD1650EDFDAC8C40C1AED61A37E9F6BB385C0DD1D00E5BEE20DAB665848A65F78A5D35696F26FC72EA4781D678095B5C5057A716DD56DBC51BA94C705CFC053B51D4BC652CD8F66B337023FADA247F2'
				pk:        '78A5D35696F26FC72EA4781D678095B5C5057A716DD56DBC51BA94C705CFC053B51D4BC652CD8F66B337023FADA247F2'
				message:   '24F7DFB558EF7F152490099790AB1E459104F5EE6C0F6D6543839F0EB43BE582B5D939091AF67C28EF1186F6E1BBBB26E69E0D3AC12E585D00FAACD5176E27AA87EA524BD104E49F3FB71CC46C6D5FEF58B77DDBE66D6D07250B0DFF95BBDF0BD6F26441AA14DD647AF4A82F367D690EF94190F77AFD9DEC2BFD5FAF685F94E7E65242D67C5931E9AEF8D98459990585BB765F29A2C65E18C9E19ADBFD8C5C547901C83B022485596B33BDD91666CDC6D95D3CC5B40DE8AF8E44FA01B39D1C6CD2F0EB2660DEE2F73C13378B75ED5DC3E34E791AF82E446428291AE51BC16CA3BF33C6742AB015527734F3F87111D8A82A16C32040DB9F986515D775315A2C2F0CA89C4E9687DAA66EB9F598C7AA7AFF9F4B3F47F1794B5B815DFC0456830C6DCDBBA3EB1177F4695EB4998C3721F6611A2DF93DC7F9EBAF94ADC68AF1385A08452DBABD0B942D98890641DC29DF0948E8ED3CB18B519A8779AE803E107D6F9F91C26C416ADE4F57DF848F6281655E14ECD60860D7ECCAB16F249C5BEB0C1C1868C24287F4F61FF04E149E560309AC15096C4B2C96D862D34A603789CF9D6C7DDB936C2E7A688038039F393AC01512A6AE6BF8588AF7ACD5F0BCEF742E2290884F5E6B16B05A8102C4D52442AE539039D566AC5F26BBDB46A91D88FB6A440D28E2E78D504EE70D5ACA1E13653E55F279B85AB93B4A726FDCAFBAFDBEB54B21D73B6398A0CD49948EA2F6D295978A01A7DB3D478C1C488B7A885A9AE376AF519CB4ABF040FDCEB700E6D584D6EDF837499D736E06E8D6822BA3956F844A7A6426CDBF8ECFD49F1B494430629E732F10F7DFE45EDAD61E5C437AC5DF1818FB314974F805FDF0162EFB4E44244519FCF083AD87807BC4D81ED3BD7EE5039A698E69757C9B64B2BE7F5F6022B3F5F119C15FC87A81A764A7C5105CB8BC6F758F1E013A165FDB5CB9FD2F2EE4238AE97B8B79ED5A93B96BC87FD557F81DAFEDAD4484AC9C707D93AFBA5B33EC6FE47C1D087A68A91DB914CB9EAA93F28A1615301C9EC9A0A8F2F5F3230A14A784097313C7E20F32E00A4C0D24558E6670B7BACE03B7F6E3F8440017AD48B369C738202D1104A945E518E81281C1E4A809A33CD773DBDFA43785177127F44BC91CCDCE08FD980AAC8E2EAAE35C2D680FB5280CF812D03695411EC61BB0387390FB4540EAD19AD0169B4EA8AA7121C2FDA0C7AA9B85460F5DB79FA3CEAFA5FA37D91B041F2A09D760C3913F212EEE35E4EC75C1AB704CABFF646BF3A8FA93A8DB6FD699A705AF7262731AE7314673C8AB489D6257816A0E72C20ACE9C6C4A7AAAC28695F69A7E824ECC43157EBF6E0933075FF3753E6A6104CC332587FD3EA58898A69F50A7D00B3B12A0C2E36FDAA5E891CBDB11D3135162D73CC6A5B995EF8E26855965579BFFE371C68990CD394193D8DF1CECCDCC0DF20BF6ECA6B37D029C318F1CB06E7EC7AEB8A8DEE1055D59C4E27922BC31201D4335C7E31E4AB78B50A88FEE26FD230CFB9B4E0CEB0F43B9EF15375D3ECDAA2B1FB61AD47B7A63FCC593EE24BF4D6FFB40B8F0675C3FD45D09425E81477C1F3ECD4E3B95F863C5EB02AA4CBF6D4DFC4E977EDA5E0C77795A4C1237406666A711525B72BB9B067A1A16FCDED59A20704183C5E7EE8E72993F09D79C727EDCE8E180E6DFDD8F7F137F6D68D0A6B68331E885B61D4E4727F83238013AAF85E783E7A29559CB08F5F7A0132F1586A4D2404486225A01C48A77D9B2E8D3871F27AE83EF7578F7C8B70AE0B7E1D9BE00AB1B0C885AD6346A725C1B8D218313D6AF81ECED1632BFDFC99E5C56C57421A504FA36FCA936A0149C99213558C1671361A52B027EC3FBE117B5BFFBEAD0049492734F8897757BDA836BB11113D795899A4627C908B3195383CD712411247F4DAB340CED4A015A896E34B598167EAE89DAD01F691EAFC99E619989F1FEEA0F3904C790C1606F59B9B04678D2517AED0DBE700E205D83153BF66C5DA4BB0ACFE7060612038C6DF9E9F07DED34EBC00ABE3D45FBCDD1153F16CB1C2F59594A379E7A63925C392B52BA3DE0359D9AE15825C6B6EEF2A8494A99634B2EDE2737C9261B881543E6D1752C37A3171CAEA262FAFB5690237152278FA7782DAE578A5E55FCE440FDDB547C56D96045CFD9F21290FA8669868CC50B5B86F19863274F8C7D73F00EC1335D8164DC1CE87CAEAD803FDC55FDE407D1460AA5735A5DB95973C2DDF37D5A32EEE5F76B7057D2D0B1CFE14E51BD9B126971F04B40AF1855ECD534EFB92E7D8FCF9199F00F4E78C2914B558CB0498E8E627C0B710C29C387D607B9E919631C065B9197E04BFE8E75E2FD740436EE5CA6BF4E52D534D9216671E4EF9EC45BBF06508C7B0CEF4DDDB552404B2D90356CC5A57D44D9696C92D79E872E28B3E0B62D2B0539A3B402230428BC42C7B0BFEE9F0DA27F7A89EA0B892F2F0F135105719508FCED7ED47A6825F7CEC375F6C206AD9B802E2575BE2A18840E1D1C271BD2EC31398AB76D891F3CC7F538B3038F984D4B362F24F1A2CE92B35A08F4B62F1A3081C7048F0F51E4CAA41FC74450DD738C02D44C414C54B335C89A095154C45C8F398990761B9B2197787B78A4D8962CBCAB5CB812BF53B9123D202A31E95C461DC4A0DA7D991FE9BBE70C950567F156F2CBF2AD9BE1203013062A96055708A30D81E0952E89F8AF59F89A33F067C03DD325813A8D69C8FD5ACF63764879E1551AFCFCC6A4C57B7406801763DF7AFF777D730FE6AD22A00A48845AAAFDFF2F705B79ADF0DF3DB0E30C2E5D2D731082B579617577E93DCFC7ECDB0455A888A364AD8B74612F79D9F2EBF9247CEA8CE64CDA0232A063DCFCCFDADD6AB8309CDC30AB48BA595D5CB7AC02D954E60DAAA5569435F184B84EAC67E4D1BDE726DBCB3FDF31278FE37A81CB87EBEE0F44E1A198C59094FCDBBB61D2D89DD4DF273F98F1E898C7AE426AE72931CD3F1A208405B9B0E526BFCCB4D8A6DF69FACBA3B398C6060F944A9A527DEB5061B1B461413CD2697893C0059F007DE36101C056388AE381A05B5C576E3144A62C5ECD32BB07E02A50032E961A67626BECB9CC962318AF2EE370692266236CA629DB6C016C699C2D97E46EE7B9C6F20A7DC37ADBD86D8199603A9B5835780FBEEAE75D0D71E02F6694A404A5B10F687FC89F9A76E2568D87E8DEE19BD030D29B891FF62146BBA918395C3165F4697741D56C88081499DEE109A3C81AF869C3C50AF90E28503EEB51A7AE0FC038962AB0F9D90593F6DC9598484760320C50C7491D69FC1F1A701BDBFF7EE4A932272869D5D46BBFB3E02F061929996C1AEBD08B5842E8600000856499B87425E2AEC2E2B37A1DDCDC1F8C06CAFD209FD4B59373A4C757F40ADCE4F3B147DE3FE7FA0339C86E21AD5F7553AF36F23DE5F436AB78F75B20E6E88A50D5287C522FCFC3F908E214D6802D8BCEC5AE3F7F5AB20D700377AE02E003E64E9EEF4F382E3A01EFB54DEFF2643A2226FA3B23CD36293F2461AB8C30BE7846F8D57911A354850AE87B76A89AD66E1B90A76C7B26FBBCC8B092A3BE38237C655EE8C6617FCBCA9375621E89FED9D2C81FE3B0AD24D72FBE36F9DD6EE7FA6C070475826D9F8EFE4055905256BAF3C18D018BB8A42B81DBE05665EF7E0C2024C7B8D87CC067D454D888DB2EFFB886242677E98E0BC225E08135E941F366861C83900ADCDE19387690977ACA0B0210CA9859550528A4B4D295B795F8DE64EB5252E7300F821E7E7C7D1233C094BA98162EC7A6DEB9D903B4A08DFB5D95B589C3570F85A4193E923E380EDE2C58545F90152BAE67274262D78B494E145DB68A5B3E8B15F34BAD42DD2FCE211BB08EFEEFA258132011C84F6C03D0525B1BC10D59298FBB564301E9284BC03076AF65A8DDA56AD66A10B4EBFAE258F535D68E9D5F45D080586CA35979C223D5FDC231C5F80628E9B921522AAAE827FA9D7AAC4C20BDF2A8745DAE068E23F8BC3A5FD321DDF670E123AF5B51ED45DE0772327C717F5E34D0E30EBB68E74C981473406F88EF992C1AEC2BAB548ED6B72FC6965227386BFCAAE7C3BB09105C0DCF04EA28A575A49DC459B5DC7C091B949F18CBC5F51B9CFF9BE5E52D8C5E86CFC8A7B4702275D0FB8C8B6EC43707E28F144F1A90DF25B584740D9D75703028331EEDE45E9830E4B9A9ABEAAB9F110C395B555DB591A4BCAC064D'
				context:   '21F397364A4FFE1004AFF019B855697B3D4AF50F2E694DECFDF168A479A5C87D8AB68B13F5E90DD5484BBB00C55B35950C0A50E0BB7F70AD078D205825465BBFAFB575EEEB75868D2AB08F9F1754791D498EEBD465783300A577897B773886D7EAD2543F797E'
				hashalg:   'SHA2-256'
				signature: '2B2026C74F1F064C35DE0B08745BFA7EC60C0EE1B2A758D02EEACE0A119E6FFD96BD437DCD57487B7889EA7683D211BED1E0F7E456FB5D1EC5608FA8646D8306364E70EF7A96C61C7ADE39B66B2770A169B98982CC74E08EF91F4A12CB9ABA2F21F074061CB74F3F6725622B07C9CF8A4612A8BCAC2D8AEDB477A843ACD96105DC9E29A2F0AFEE6367805D69C65DE04581F36A6346AB820A864CB2C1450619C918762F8261E733016385B47669B9F700DE4D8079647F5576E5B0AF3A3DF5F77FA6DE7896BF1CAC50844750AF806022718BFDDD70F78F66173923DB4B0CC65ACE5904C493E6294360811EF86BCA654E5E3C7686AA065C45663A4E5FB9EE1323F148EA5153718C7794B3635879436FF456C22D036E52D6631D920AF0EF73111F54ADD9EEA49BF52669614E324942B02EECE2A816E17881AED209F57864BEE05124F32A18455F5A019F6DED258CA5A692DF58E2266C7DFA37B4E1FDF9620995AE67471D85284341BBFA162240C1874B07082BB68FAB35E0420B98E427D46FD219E632BCC81EB2D730C25BD293E0DB589BEA2FC68260DE6D8DFD706D0F89109C5DBA8F8FBAE2136919E5431219047D6DA5BB932B5A8D724F3128B18E8575E0E7873B17668F9CBBAE4BC222FC36942259AD3EC0E50D08C4041E737C0E85986F6751A4C945656B972A794F0067F3DFAB921F79624F519F3844A747DAFB77B82CD02B998B1BB710E65EF8F363BBCB7F43903561389C5AFC80624B6723A3F49E4E0D0F1AFFC072CADCD7D340821523FFDA5FC274FC23911A76E0AB3939505A49DAE63A2BA5ADF3E740EF3B9EAA4CBF6D2BCAFD4DB5B1BE79B7A7EAD82EF77E0BE2B66C0C62EBFDAF69792F71321A2225BD81E2CC1CE6FC5AF306DF5BF7FB444FBCB1F98E1581F1D4CAA5B19CC442547975DE63229FFFC4CD65964CD0FCF0217FA47281A622451CE6AB92F52C7B19462BCFB0EC45D1026E1BF18CFD49AB5D5A8C617FE247C51B90CE1DE46B4318AD68B67280BD832BC7A518C6A76E8C6F5AEE2F99565BE39179BB874303447DF78D1D4D3033AD34C025C62679C51E80A59E1BD9AA3D7CC659E8777F890E02DB5099F7E5CD9A312BADCA0E73C591B8089ABBB291BD5FD6BAAED5BCEF7EA57DCAA90DAE8024302C667354B6A1635FE0032E44B9DE942067C366651AC455DEF126606C3AB908FA051A7F815AB503D7777F27374D3F81DC535FEABE37BDD76A837E536145B1051F057873A40F24D57099DF2A952F24F037622F2B06EAC3D6C221BF6180EB1994FB127A822C560564EF455804B7E853D96C27CCCC12ECBC214F791267C69FB91B293A75725534FE3AA315F8C48DBC202E9CF8874C8F6E17AAE756BDC42072EA45BAB36EE1FC0116E7CAECD92B0818BA263E14B8C99466EF081D4BA702AC467C1D7791CC27B3B14ED0218DA9E91BF54B0F34C6930AC15493AF107308D0067750823D0CB3F87A357AD59380BFF311F49F6E05979852D7DB2415954AC374D81525B756AE1672928E2ABE2A813C73D080ED456774F47EA686CCA7984D25E05B3DB747AAB2F639C4754671B42905A409EF59D5DCC5D94784E682734A451AF4020645E58074212C0CD3F4ED161CD593664134B375475739034690466739519F1BCCB07AAE9888A03BA435FB4F701DBEF15434F716D1FAD6460A1EF2811770508ECC5357C084D6D6BF979F1ED031E71BCE114EEB02FC0BB61DEE40A5C9C1FB8DC1F171AA00F5E50B17EA705B38E3DFB67A4FDD9C5774EC7EAC07BBE609504D0D949E17BFF1C9381DB48B0B19C2BD7E021D36A5E49178E1C031A9BAE9695A05AED4FCCE937C1DC3CAB2807467ECCEDC0BC81AF7921C5E9075B48406DA0A750E8087D4C4193988F22B6D316ACEF7D2592226A776CDB93A9504A16CD0A2B61DBD032333EE4B24D9C8CFAEA2CA779C5AD16ACEA72672F576A99A57D8BEA08C0AC0622F7274ACF8E87E99B9B758CEDB3F16719B2360DF4466E33903DE94805B7503027CCE748193FFD5345FD7E99FF87075CC1A639D01444515CFBD55D08B56E4A154FA229804CC39407DFEFD263E4B61C704F921CFA3207B7C70EDA34A758DA7471A34BD40A001642A5D47A9E20F8E48C5FFE20FD13F57C7EE22FF86A574730A1478B4A03F8071F682D57E7567E49B9671FDC93B3176145F437A8637BE6F25EA39253B9AABA4D348B89193C52C1B9C368E9D55B1C7A92FD2BA564F27076851C55D46FDBB95CC2F4D9D20A95E8DD6C34E0F82A849CDA2D5C69E2D037C881B2E62CF4F36A5526A04F35D26CF696820E4AAD05267A0FA8F196CFE4511F00E3C11EA0115FCE1E636C36E1BF01287A4428C63423D38FA2273C24A00395CD233C239D4E779B3F475D7A8750B7C75A440454B839521127EB9ACF01B472C261E6B0F2C84E4D407D6B9E9A3C379CA524A29013A83D5EB8AE078BC9B519FBCBEE5052C0664536E3EEEBD9D36AEB3F3E2DEB2F6A04D0BC6AE0C9B3996513670E3655C4F706D8FD34FFC779BE44A6CB93471D53DC87FE79B611B4929AF85C9C1D5F24082A26C8815DBC43FDDF97DF7144143C84B4AAC22E2B3436B049876D8336E19C3CE882E526AEF832536DAA3704803EAD0CD59705B158E094D51892573409863D8D5CBDF18D1D5892ECA13B8E670497A8EFEF7282B26613167F64A7D85D2660BA52476A3201A5D70A6ED749D919539C888983C88DC6F43836907AA658B2976745F7AD2A0108445D6DC34FB3C7781C949BCD1E6C80D61951DF52A4BF29FFAFCB9A12CB2F3FB2E78036A790C41E3C68246167B44BEE659890D47A5D1642D6AA25F0BD68A46AD316164E65A292F9EF3A7358D1864EBA647656AD12FC81B0CB68412ABDC60DD07D1A7DFC3FDA18E6A86922EF204BBF2FF3AA364FDFDECF4661C3599C9032F50734B38B26FC2F39DFD5389116AE7288AD3EDFF00A4DC398EEE63CF74AACBFE3913C00DB8F5A2C6ADCECA6B8AFC0CD3CBD58945138A60CE3CCF151EF07E34CAC2486D74F99C18F0964623FF8D1705B0380953808FFA29793EC9E4DB05F43992C271164DD8B4E4E4DD7F6ECEA9526F7D334003AAF18FBAEA8A35149E291D513571FB01A5AD70A63FB6DC983718F307D9D311CBB9F59088F1D0F2104C6C5A65AFD36B730F7B417A0F4DA00DB1E3A1774CD1FD58D02FEC00B4BB2D4038E6FB6EFFD830F60B0F003309878ECC4D9F5F34FD3ED34FFBFB4579F1D672404629EACA81D7318E262D517F926C3CECEEC1DCC0B0BA8ECD5AC4385E4D48BCDBF130957F50A68590B6AA450E5BC1817B3ECA6777E7BD1B2ADBD3C0F4CAB25438F1E18802F5A11B8D07B2D701107FB8C44FFC5EEE1D4B8F5136454EF4702CFF706FFA33EBB69719B2F9E454DB0651441C372FC6FB461326AFC0D645E10B8D6F04B033099E587721B55B438FDDC6638D89AE387829F027D9443A7587CABEA37E611ADB5F63F4B960D86BB675A5316304A8C1FCA1A6C108A7C63DD09A83A68392383AD90840106170B5326649380BEA58AE3775443D9D49FAEC6DC930F7E0E1B2D1FF3D987686EF7572247CAD7598E26B755CE6713D16AF14A09D1AB9197C51230DA39F83C7700854CFBDFA341DAAEF17EF4D1314A8EB6141D0E1A4225071AC8D89E3873A5924AE746A9AEA3D3A60F129BF6BB1817C50CEE01C6789B8612F5095C77D405A5B891FDB32135E63C98E592CCF286209E380C61802ED9F32C89C321C211A046B950A694A29AB5A113FF59CF2483C8539186ED406EB7A977530E750B90C4267879874F7E1683C54B026D55178B9D3A6458A3CF2B7F709426E02A2DA5A1A434626F32A67159D9058E3FF8D259B97E7439DC74FDD6D06D222FB65BD611125605B726A2EE97071D61B35FEE9AF6C7592D19ABFFAE7068BB6FD78BA4E27A2C287D81C1DFE7E189C15E3A612802BDA054854F574FEDF3AB9DD87B30268CA1042CE0C5A404642D717AD27A4DE011E97E65210619F73878B5F770C1BEF45630C767316D09925F622E303F872F0FD07742297C4A41F8057E6E80B4C11DD46752E86C7FFBF6C7D81B903ECDFCC1C2A1F15B6EC25007A50A90F4DCDA07468C009E09410C367B31E6F75A38F30BAF10A51B2C87171011093FBAA18F57B693586FAC79702CEAD640C47BF055E2D4F819DD2BC9004F364CC1864C8F0C9397EEC89161FE1F4DA5EA78804E97372176AF0433F55A204BBB1AC08C1A844C0FF61445E5257F38CB3227E3D6742B24BD11ABCB406839588839AA3563E180743897DD05713D06D7795E33B514E0870A90C976D72565028A7BEAB0A6126057E255F9AE197356F7386E157B4AE52B8CF4C7A14598F6627DB90DCBE634C620D77FDBC9A2548281A57A3FD3FA6A49ED1D57CA0AB37D30FFB7C9ABA0C1982F7D08AC7ACCB22878F9D9A3A405F9BC3689AF9CA431B06AC9866054882439EF7F4525324C06331FBEAF71441BAA15F1246D6363788CDA2EEFEE623ACF1FB5643C04A3061F218D39095E082C01C20F2765EC21BD9D25F377B143B6FB54A353DC7574565E54B7E0BE4F2E061C473EAC0A2AD9FD33934AF48CE71AB6E9D4E8131AADC31E95C2760530A74E2C1C1B0D24303004517B55BB186A65506D2006CAEA93474AE7A2CDF793027049B8B063EB359F3F31C8ADD9F4D562FC9917554566903F63D155DCE937A306CC7F2CD37FEA9EFFD260BB58632AE18BD40999289CD3E1FC6B568FAA4E8B625C982F52EB62030A5A31AA3332EF7E12D4E3318EE3A1CA3C03D12664FD6CF53B17CDBA056D244901DEB2585DEFD8EE9C8BFC7295FE0671F931E55E20A6B96E0DA0965E43587F0040F66A2F4C5767C289AA61BCE2C839801C23081044347F595E0959F2127EC0B0B6600BCC55B8BFBDBDCD70AEE4F1AC628705FBBF35CF09671263F5C787CC7E95DF355DE629BCDD8CC3933627BC3681CA94D569257B0A823AB41619D65B4EECBC0201839FBF59FA26510CA150676D089495E1890EFB97EF1448A7A62192156784BFD92D73982777094ABB781A9CEA8DB0ECA84ED82381EE68C456C7BF44ED9B2CDF141A8C06AF9D23101554C8CAFEBBA286CCDAA5B138E43967BE5037F41B4F0163EEEA48802506A1FB5FDD32997BC9075D23CF9E4585BDE6914CB618F193393E01E793FEC71A7C776E364437865DFF22F1A85BB02F7D6C03579D9729BC50C2084ABC0FB7633B489984162FCA0ED6DCAFB7FCDB081743AC7F4617BA8E1FDC723230956342FAA591D508C5F325542A7B77E231EC5F4B63D79EF0540851D6D7C15DE1ADBD873593A664F4FB376846BA90565F37D4D8533FB15E4874816A7B61461D1F44DACAFB1E9755DCACA1E22567DE205CF41E7DDEED4D1C8CE0C4EF202276A42E23048B0F5D5682B54B593B8CB65CFE511F2DB95D7E1CA64A3FF4355058CC3118793EA8E3FBBA72D292AE70DE4BB17F730BCFAB8B89259063F2CABC46EF0BF57BC7888E0F152D208BDD44A0788900DB8DE575E4CD4D29CD0D23B31ACEE0AFF0CC52B6E91F3F38AFC5775700FF08252778B1AFC41C81A86BA74E5821DB5169842D59C0B20507CF48FE769AE8872B11EF298FB80FEB7F70D5296A97666DB129A5E1C63CDFAA664241C90EFE73CBBBA48E762846FD0442400519B579E79DF9D4B7CA9CCD241FBFD1318A1A06CCC88744DA254E3D25D3663C75C5F057EC2F8877C3EE2EE247BCF804C44C5D110DF8F8B506834FB1033374139CA0E00B63DE7A883A27D67393834167FCDDA5EB5BA1C116D6D9FF51E55AABA47B4A885FBC213714D6B20878F8788A91BBEAF29968BAE00522E4154223AE49A88EAFFF53EA719196EDAA6AA425935CEEDD99E244990B47309B2975D76F0F48F1F68CC26EFE59B9A49905F4A5723D1E9607E3019C4BB1C0A437FDA480C4271350EEBC53DC6D1FF793FE96623766294B58E270533888FB672C970107FD1AB2D6690E792E468DFECF1A02956C433FE63D1FC8497154EEEDAB685C23521F2FCE8CBC6BCFF157A7857A03E50E46998E3BEAD49D6FC8ECB0C9381E0F66E41B52C8C6BA973E7901FB369E8CB17F3049066360D21150BDA5D2FD95FEEC9BCFE7060CD0A118D8748EABA06A49D0982FDC8D91FFFAE90C1747A16A79BEAC2621CEC072B62136DC7636868851DF267C3E6A2416DEC090ED6B3A0A533C8DB9103F88485AEAB1C44CE8A0526D097485ECFA7ABB10E0CB7698873927C4A5C0C7873B96D3D7CE190E5DD29F28C9377EC8A75D9516268ADF592FB7AD139719C6C2147091677DBBA9C4508F619A88271806829B618952BA36220824F967B7C82934EFB17C193FCDBF9825B75E11EDCA6FC0CF957ACD53EFBB2648CC33548BE49BAB6F7DEAC34DD474D17ADD9307F2DC6B25C57406E835CA291DC69B9BB8909BA69E0208C68B228355E0C83130CDE33C4A70615FA014568A914143FFAD6756302F85AA87D7EA07C536DA2FE7433D02773AA9329F1E585218723071DDA196F08CF504AB7A7D9B674F04EAC1603EC10C0AD3D21846161336F766AE09E00719080F2777DDB6CD99023F504FD867D151E376DC60FEEE8F614457054B72596418A935919924E1B381B7F07554FC0EF7883546A2D086AC549D513E391CD0972A41B890EB5A6467C25C5AA836EA985679A25E1D166E0692CB69986318627059C879141D746F8C19C0878A414612DE9AF8CE8876E5759E6ACF34B7A73C95889FAFEC24C6CE6FE9DBBCEDD7D15F1331682C43DB451AC0E9B7BB48323CAA77A5A0036EE3F44A0CA994A6335884B426B51CE13BEBF53E4739D877A0F0517AD918D902121A630709800C2CD0133DECA282D194FC38249C36DFE6C032E84F19BE5FCB06C8A4CEBB4A2220C9A7C3B6F34A08E835C64EC36CE6B216FA265F84088D4D3B191962594D6D34C066160FB0AD2FBC1534068530C8749CE155AD45ADB453C8C4E578DB31B41689DED46896EB39FC6DE9160592B476B24880BD773BBA7F352E51E8B47A463B14CB093F0E434277B499BACF4169BDEF680C3C02902C300530EDC39D69013C7F6BFE068656742511F13B0F2B8B613CC507C269D725475EDD2BCE8E530538A718AE0420C76DD2BD6D62DD076AAABD78E6CDC8796115D1D9A384E9DAE11FEF21394239FBB02A4E88FFBCC8BBD4DBB00DD6B053EC073944336E989CB8AAE1E338E38D7D8090E0AB9BA1C2ABFD1C8815BFC5B18ACBB89264D5BAD028B8E0E85BA1D7179D719360360A87901C1B564C1345264706DF0189AE1F140EF411A9060A52283367EAB647B497ED4BDA437E495EC17B7F9ABAFA3E0C309128652EC18D7949B201904B566E156C50E17932EF4BBF128683BE3DD52A946005A14EEF1D622524866E69D45D96DB51884085D0C676A29F72CE29EA6DC8FC08D7F8D746B026318E8E678AF1DA04796A3B4EAC8BC2CF466002CA6CA4DA67CC125513FFD06F32524281B740EF886624A5E466FE67BE817F266A03DD32E66752243CFE0420DEED22290A9DC15C59826688D0E1AB99E98D2329AB0DFEDA0825E025839214E1044158C844A8C4628B196B2D4160F0A0D8330C067743F657679A18A8AED2EA7779A6B43F248A2D9613923E33C698EFE0A555546C38139FF95DC0EA855B9B7005CCBE4F95528B594357D3A83343572A68C4F3A5F6F2DF91E648C10BB53B193E8C156DEF087BC9B38645430C219288F41E8CA7A196B6F3561E7880496B249976544896AA7B84DE468FBA51FD05705619BBC6BAA943D7A87DF382F40E9D1577679EAF1CA73136E6FA07E5EEA8D3EB5F2D99735BDAB0C4F3BDCE9CC6F6F36D46D528B3E44AE71B78E087FE4514FE8CB7B57EFFB5BCB926DC7BF8ED74462C9C7280BBAB6740C7485BBB8A5147A33B22F76CF026AC9C577BD6D3D34F8ED69D7507AC7A6DA9C159BEE62DD8B5CCF069275DAF83EAE5E43DFEF284DFE96602508BE070A91AC5FF64BC2A7F35640F540DDE42D2AD4F6A5B77AAB0770D3AC81EFC814ABD15C3888213D8FB98067D45D11382EF6BCAB523245C4BEA42DB42468B0324A383E24117B815C09B1BE08BB9B7EF2070ADB5BA6EB0D4A058F3B485AA74CB5CBE557308C591D5F5D164F61CA80221BF0F4C2715A1AC59BC2D10AE123241781C4618E5993022353C2101EBB2EDAA211BE911F270FD0229CD720625368E278DA6C8DDBD3FD40B859D7E3F5FB67ED8371AF8D834ED4C97F2F7C0C05EB37EB10932AF88663AB52CF80C5979C1123CA3ED56EA32D0B34FC7D0E6B4610DD910A2887D0C249BEE253C528534B1B994FC8B389B631047439951F9E5C0ECDC982DD4E04AC9F27C5CBBE61CA982762A3F9D08CF7787777E4EE71B803D3A5FBAE3B154017B3B7A861532A6459B9F900614DB0AD41A7C9F4C407C77DBDFEC1A837F4D5C142EAF86BEAAAF3050528B0E4AD9697D510968FA1E2FD0B90CE49AA52B5019DAB78CAA4EF121A6ED49B660427E05F458B8F036A19DA3115ECD83F59BF73E3EF1EE9A29BF86B9C6394178A165C607C7FD4AF1C815365B14965099D5F51D2FB19C4B9C7C371A55FD9A71C582F968A4A4DB1A46ACAC53F91E16976B576E7245257D42112A23ABE392722860210BBB774CADC152C68F0E146B1589A979C752CA51AA32B6DBF5B40A92377EE36D13CE3EA53593A3943839FE33F6FD0CE41479D389B1A04DDDF83D18E1E0EE8C77BAE6E4261099800DEA012273A950E8ECA1D9E084E07F910CCF0E98643DFB3F66F98427C44C3B952A7A3F43A0572FA2F4BA59669FF889C1694530FA33BA7F8DF923A5E680D7F86ACBDBFB952A15A7760BA4A441F860C50047EEC23D164C23321F851A2BD248D1C441C6DDB8949973BEC6C453CAE0D97872B8176DCDDA9280597DBBFAA1053C153E2C3EDE7C6557902956DFF08221EEDCFFDFAD8E07C6033F9877AB99D735ABB1E45555B8DD34953CCB5AD0E2FCDBC3F9CA1182C4D9684611BD9D8BABE670CD93BD9DD23C3038B1C55A242CAB5A6FC9F9239E1A59C1EC5D73F262029435E3FB47CA3A627046DF7910B984504C2BAE04A9699810275DC62D7B924FD865467DE18A3298DF5DA92084AEFED9B1422ECC88EFD648748487F2E17DB0F90C27882539213863717121A52892AF463C747626C0227E326265547B82971FD751C7AC1ED858B79FDBDAC742D978F3FD7A7B53102FB5568643783AAC5E799E57573E3D6E73095D65936728F88C3C811228ACAD050116F264C9592A8B412F07AC7AB81969D6915CEEA26E16601708C40B9C1AB0E82FB9914845C43D77EEB1D61F8C109AF69A96F60DDEAC9439112FB3BC5EE6E1F0DFAC531FAA8C02371FDF1C38F2DB4792BE16B246013AC9CEF40AF063B222A04864A49ED51C65A28A0F7DE4C316A1E332523BE56E7B02278887EB66A5F0BF9DF1F31F50D638558B4C1179AFCC9F7B3E690EF7D9DD2A815C7DF361A0FE86F9D3AD2F50D7A8AEC0C82906CD7668455C41530C5E0DD5764CF201843EA80F240831778122229BE86CC7A4BC9A708020F6EAB4A7BC15A111221EEA5372B0F4FDA307BA1275CB3FC18E18B9011EF91708B888E571B0D6E38A249CADCCC65E26CD5B43EB1FCAFF9DE67AD4C7F0CDDCA46BFC013D1F352FAF3F888C8F29A51EA2BA3973B8E7E5E2FF0E24A05CB98EBE9C9BC4BFEF6A7D70CC5D180F4A2278149654174B3127EEAF78E8BDCCFA4CC2CC76FCCF53210DF29EA15EC8F305D9247019DE35A2D78EC7392E545ACA75A301873A400D2EA3A6832A1B84FC2C29B6060C545907EB6CF3B7F4E74C52DF10C9372AC30EC781838C877DF2154E7610301E58C10573A2270A908C11156D2D5153D971EBA61840BE9FFB480EA29675157A305841E3DA2B628BDED01F4CEBA9153639EE732078C0A0A6AFA29695624FA7D60189922A005F322CFD97E84775C8574567A707C02A4826A6355555F592F609F8DDCB5442E05248269D3A9A3F6E9F6895E683CC9E3C7E71AA4C3D39D7FD44ADC23184031F460BD2B5DCC2251A145C7EAC17AE8096965F23FFC8CFA20D724087E375632F8690EFDAE7EB66366CABCB4493189293378A91D5B98DD99118E109BE7E50FB7D89F4DA144CEE291A3F0C9259AA006CF4ED8EEA5B4BAE5E8B610E56CADBFC7DB8933550B9D61CACF0951C15F302A09885BDA7E3C33EB5394C294488B4025DB61194FB011F576B3632090465A8F5173DD3F566BB8B564B8F623AE41503481B24AC7F144A18A46BA81039F5C748DB66D80A3519B4C94A203367B9C2D867FC2308C0F29AEB94A7F8C88FF8AC76BB148C01A76E0E3558012345CEC41E30176F762E56D466C09442E03465358289C2ABE99A61EE963BBCABEEB2CEA9C704E87134A7C76E7D8368C013D940937F9E1378B7E00A8D8D7268D91EBB1AEF2CA96EBC38F105AFF9065BEFAD7D0B1B6990B64C039C26F8641159F49E7C619078C3AF400DA8D54A091999CC7E8436BB93E5097437D76303A4AB8ED473A44BA5B51D5CA77726FAC862606C183D2B48CD5026CFB9752F50AB49D0D52DE282151CF9CACB3A7C24BCB7B963047D78586900B6AA181F8141A00D518E88BC06CDCD09520F28A6E21D51C601D1C8F1911C9B65DE63F00E9684A922EC3554D8B761CFFC5EA5181B7DEA031D77E39EB43DB47CDE9FFC7DBCDC20B47CEE29F62A87B4AEE2697340FC86BB61B98259A7272E013FD2A837274641D34619BDC03917C766DE4F355F54A4526AB09823547D48F9F5C20548FC71B7C40F00C499651FEEFCDB68F35022CA59F182974F57168CFD8D65419FB79A894305873C504BAF397938C6B0176250DACF808FFD2C5772972D771BE9C7FA9F3348B67323DD592DE7E2E330F8DB28D09B33991446A273A7FA961ECF33CD6B972F27A9DEB3664698BEE149F882109EE18BFD5534CB090D670111FA4A9A4164B058939F06A04ECED2B63754EA2E10F36A99543739138D2CF3F3E72B32B71BB5CF26C86F385DD4D004B790EB9BD65BD4D326E820B16765AE7486DDFB7C87936FFC89C2B91E98E22CBCBC02A4F92FD890039F72F3B0EF80D81167D4469E4653E4D51A2D7B90E7455ACED2573E536AC9001396F4015952819249386B04CFB8CB389C6584D8EF6AF87C133617D432D1216580BB59C9D40564CDAF71BFDBA08973E303535448860207E0859D4103FCD965B6A202DB2B9878C215D122A020C94F6AE051B2F6ABF2FA1855131FC33F72F26F93C81DC2472D7EE37263EFCEBCABBCCF28C060BBD9D80861534ED00E3679A678D655EF15E50120E526EA623F56802F4930E20179EF674E5CE28737E8CCCBE7F100B8097925B024A53741B880AD6C611D2C32D6C0D5F3CF2074A4AA96FD0BB1911815EA5BDF0EF464F9D0DACF5704DB7516CC30E572267D263011E38A996D631C42B3B199025AB27B424D2831688596735AFE0CE11157A0E92AEAB7C29A7F8302A50D78DA06D7B7EE6602517A9DEDB84C9C3797F86D1E20C1910B471EDA7AAEC0A159124028105A6DB7280CC8BB29090444802E456A2FEC940FBF50932CAE172B414DD930A57B9A67CBBCDFDB25FEEE95EA251C379B662055EFBD3C09B649969A45A51AEBCEA59A575BFD0ED570C7707D9B007C87C426FDF2946A2BACB7F8990647FEA3407A6962A88A9781A83FD456F6586ACD9F58857C48F16E27D0E9CA1D3462B817FD1FC5C5DC1D5566DA6A4FB261013A19BA6C642739FBF3DF8F59E7F3BDB5E6E35ACA0369E86719186D9DFCA86F056D15903259BA84B56D1F1BEE6E118BCF546A4B2E98EE48D2646937C6FF871445FCEFAD37D50BFC75F91FE18D2239CAB5832779F17111DA3F2B0141C4D0FFAE9275405AA6A2F2429AD64870DAE387E54EE37B7EB737F59D58CEFBCBC23C6DEE27FF594F33D23A58A02CFF22D1E27765A0E320BC902E4C8D2DA1A6C9E231DC4881ADDA2B3C2B9F35AED65FE50CC3175CEC55A637459D64AE1A1EB4DDFF3B5E925E43D5C7FF2EC4D13CDB71C0BE26FD8DFCE0749AB2016B09A5DE9EDD33DADF27C32528E3B48F451606A3D7103BA7007AC22A7973571142514BD8AC71EC6554C7CD8C34A3D36A1D5BF0515B2D1BC4C9C1FB6FC56124BAA81EF7AAC7B18C7FB7303CA66C261FEDE481189BCA0EF3E97D72E53A4B1EB47C8B8B6DDE38138DD8070A2CE58C3DE28467EF62178B13191276EC0AFFBF5D8388D72952E601D52C091BD42D507AB2AA6BB2B36CC3BFB2334780E504B340D61A8F3B3A5C609A2BE3CD097E836CEB262E51BBE334C4FD32C0165ECB4B3D2F103AA36053DEF00444F5B0E764D0D117E2419B4EBE0924852B36740339B425BAEF326F7638CC220CADB79BA4314F49DE99BD45FB189489CEA005A3024BD9DC022741EAF0CE0437E675415769337393D35536903A1C27EEDCBB27FE02C73AF10E6FDDA848243044D1BD2D161EADD6912B998EF8207697944CD984F9CCE19D857B7D3D7C5D27B77DD81833D6C9D32A5A6830C77A145DAE66D63F8D1DB4E663D93833A053976A0F56FA73E060FD0D575920A0CFA44B99472DF58A662EF305B5118ACD5E59D879F225B5ECB5E03FC8420812522F84C907DE6A6FA7536C42F4CA7D093E1BB5E860144B76B51905F83648002A0B6F80FDBD97244ECB0393BC4BD539EB486F3543D532572B51A092A56639124DDC899E837DA607F98F44127AE2CE58911EB4F5A22B4546FAE97992D1553C6C0BBE84F595D5AF6FDBE7DCE222804593D3614B67C9EAE2AD38C25669720F24357FA555CB55C2C72F59E89A21772B12A4382A1A45F653E7954AFDE383751ACA96B12F9A5226F21B3782DF15EEF6FFDFC104A821182ACDA277E213A45DF7C789A7B83C994C97AA59022AA5074C74627D02AFF75FB143AA6631FF3C0EEAE59B4865BABBBE6E9ED3FF4A1D81FD9FFA4B7555BF39C69C2DD93A63F07722E9C56E3452F7E022BD63BC82AD4DD0C9F688D1656FAC245B30EE7CF1AF075469BA0DB13354020CE014AF245DD5B2541DE669B12E01F30E0FCBF206BCEFC88BAB92B3BB4DA5465B4CBD4EDCF81FC477C0F578653D8FABA43A8C9F387E6ABE093CBC3848A3E166175AB2740D2CB38B77BD10D7B01ECA5A8C3F2DF39A9088E0073FA48F5AF7455131F8155D78381B1B12F5797FABF457ABE63A15CCCF0E91871CEAC83F66ECEB3A37BFB546A77350459C49E01518AABB6010D3CFC8664983C9F04256C95F297D3ED44D5F3363DE3CC3B4096D89B972146BE7C0D88C830B44F88FB9ACF668AD6D357EBE33DC3CA6B4E9551764CAB3C56885A024BC650B53B3B082BEFE54556FFC0595594E225C7E7DAE34D1C097AB06FA1EE5CB4CF3F00CA9141BF13EEDFA3D36D0DBF515506800DDC6D80FB271A639176B891877106B57019422E37F9AE86F1080600B585D5348A2148AAAFB5B285A99096A5B4BC85582D7499DA1A65AE2D96A64539BC42B33D9303E0846FBFA8B623A337C2BA05EDA8928818A2609AF58B47311298423B60657C563CAFBA6D2A843C8A0923660E135080949D8FC186ADFA7C113185B31B5747FC324951DBE69B0B8F0ABE4DED7AAC10CD7D9CC7418C109D4ADBCDEC71294A193CE13088ACA58F43928F8DE3F6CF3A6F8B0F925FBB38CB0BC6288E7FFB790CF67F02E73D6F73C11241CE24A0C456CC04429B4EF29BDD76E0EA69539CBDE79CE725F1E484B3FA14F6C0E649ACA983A05C1B55E4F78726C7BEC2636165D7F89099EE349983905F9CB1009476DECC97FE598D4DB9E06A2213A656DE00DBA57CA808293284412786FF35F1DC9DF194812C712E6FB59EC684077984FCA980CE319E3A799420543984CEBBE1E020BDC6E313F3EA602C0A4FFDED2478292260B9042EBBF53195512BF068FD1B4A8A65689107A6373A0BE82E6DEDA7A063C1C6ED4DB9FE46D48548E35E2D986022EAA4DE38BB22ACD57F0B127636E316C581F7BF7A3B60B3B3AA872EE9082A8A0C675477B83E53C9388B7830FD3A11262ACA6DBA272B8A6AB94CD6B4FD4CD7D8D6EE7C9FC67AEF35F33441215B9E87476A8D08F22DEBF6C70CB9C34722B18CBEE8DDF8124E1E3BC27E6EA2125CB050DB1D89FDD68A9C3F39C0D3F46D1B2B7A58907D6BDC7800B9DF1E9F6BE45F15773CB529BA39D8F18E953D144A4A0455FE4F6B0D607EBA4045649127ACCFED5442012587F1E0A1C6DAB40AB3F53D3BEC712F3A9EBDFCC583AE984C85F98A81DA55A6BF23190F2FF6810A656C58073FEC93329953A7842E00216CE657793D17E0EC3286E6876BC9E0611C8BBC1019F984ABFF063B85A400902BC012DE369702470900DD2B6599DEA89B28397E1317A82358087212AFEC3AA92B2D9549471850A9D5A4A2624CDAC9800D60C48A4B73DF2B7A95FB5E17EECF432CE0560EF23EC5F41FC558164D99F2F87C46576FC8210FC8034B4D9818B0290983F6419F9053FE6A9BF64CCE7492CCA164FA735B95A2B2BDB1D072F3852B1C12C9CBF24C6E6EE304B58BF1F96DC71FDABED1368FA26DE8856DA76F29BC1573A0B0C624B624C6AD1DC9E958FAD02658F9A80C0077AEAC2F15E72D67ED209989BD5CAB47DD2FEEE5F9F6F5B8BF556736BF08FA7517D880CB928A41E67DE7F05B450AAAF3B7AC77D727D9C4B3CF4C5E7C71F39B96FC3FDDFBC227F7AFB9EF9F368EC81C96A02B5567BAABA5D627D3F13E664B64FF43F112BEA05823CFF8CAF45AFA44E8F208A45828DBC31DCAADBCB9ADABA301D32A5F125588E585C460FAEF57860865B8F7AD9B1A69550042C0C310567E69F2727E39A7E10792EF78021C2E4B314B0316AC43444A2B5723A337E6D5FBB07218AA1156E083F2ADE6A1D4A129CDE035F8C7CDFE8F65A0F20377A1A2A2FD23AFD878EC5DD819977364C5478F1057CDACBD49154F940DA4E9695AB5E1F9346366856CE7A410975CADCCA7FFBD439D2125F8C99CDF96174CF4CF93AD7136144AC064B8646E87D2D9300D9126E07D4B75F5DBC2F0AC440A88A595CF428AE513E11DCAD27C8E371B682F3F7A186C775C96331D177552220D617A2CB4DA265A1359281A2DC756518D3BA5A5DA0BA948415D7E8003420F82CE47C3D198AA550E3268FE7CB0BF06CA5A421EF7DA7E88A505EAA7B387969A6B30BBEFFD2C31D531C13A7B7E6F981CA82C70C33B8E600E2786D418FCC3AAF39B97D775B50B8E2A8B10D7F797982FC80A37DE63B7609343F82E2BFF3404463FE02987ADCCC7C263B065F13F7136A43CA243FBB75751B62AD8D3803EDF8D95D4B714E3C153476562893FF80621AA2F798087E0329EC4186E4844D64B23AE465DD12D812EBB8981100F0781C96C057A3D7C238A14402D40A9E6F178EB1FCFA893AF64AE29B213E46B75805333877F4A0A6E560F517F92D8C7270F7386B848C0BF2FAA966C4480C3570F2CA70CF0116044B4F1BA5AE6A4163195DA44320A7980C607A252DA6E4C32524A4111FAA0F63EEBCB3BE2E7BEADC0B504F86E7B3AE87B1F2640353FB88CE0CC0B66005AC6C7A595D09AF39ECFE82A9E7E74D58B25A102B07D1E5205ADDDC9523BF3A766D582A58EC79D38F23B2E838B884B637E342CC630D2F44BFFBB4502FA20C43E58D2ED5C76557E782C1727ABAB50551973796B9B5F2F78F6E598CF3B62A860654D865B19323B953CC8623E3D9A334086C8EDC07CE758783FD00390BDB5788AF969F01151C368011BDDA882073B1B07CE60C99499C3E4B323BEF7CFD0BB62E82510EC99347D187F9245B518EABCABA431B9DE5860CF4554B86EEE462948A9E833D634B99A6679F0A6418B14D8C1FC642D2EA331B75D855E249B9C5DED23FBF8F5B7F3A7D3F4DD98E69779FC4BFF7A0F9ED736E1FEB6D83927B70A45D7659E8D2858658C50D43FB5ECDE1648505FF88A8A16924B056CB9BA2DCE0B6AAB71FA94ABD2EA078830D79752A0AAAE41F3B62F65D00E125FED62723E19D6AC5F07B4AF3BC98A406146F5B7B6D014B2CDA1C0AFC16F8D919383E5575106D889207E114558E8CB7CA4CD4779109967BFD513F12F18F1576880A0AAF1087345C77EF7754122EA009BF60433C88EA83864024AF7F40ADEDF198C116F615B68FDDEAFB15C088D20DA70764EE530117735B2CB37A32C58E198C3373C79F31227B76DFAFC948A8430F284FD38093FFBB3CD5DBECBDDDD34B8CF54EDE25E450EF8F5DC956E5EDD92ABFD274DE83A252ADB14B5D83ED8E954B3D9EA5B96CDB07520EE7829AC5DE552766B7D1878A3B02812C5C37DD5D1CD5AF53987506A7ECC406E36BEA257D0A02A224A5A0A1A3D9F1F648B2D67C021E33137131CD9237D778A337CD75A420FFE3279B4E17A7C2E5D660B1AAD0B157E74BCADF78E77AC846F09F41F9EC52B3CEEA9AFD09C9FA53017F849B7FCD447891E0570A907C66DFDEE051D50D1A800D50383DCFFBB13B751149196D513574EFCA2D49213205D447F8586639E084995C08908AB8A05F5A480DB1E0CA698508F536CA2BD9CF5EB61DF2DEFD984168C26A01D5D1709FDF2ACFF05D6BBC78BFB536E63C556F003B66A67F676E2A84B9012D31738A64E27FF4BDD46453EBEDD4BD812B210CD7C2494E881F04EC7F0074DFA476E022BECFA39F3988A74F8A1B7B66A3FA7BE69B33CCB64B5A0E3276E619B61F6B99AA74AD65F0F66ACFA2D8074F148331AAA748124D1D7A1BFBD94808FA84D4B94151233732C08C3800DF98C22AC52F4F5863D470E6C785D47BD31164931066164BF13D2993FD1A178C7F6E6F6DA2F7DA08791CD00DCFE3D488105511F8F6C31E3961C94736089CE570A914B85D327E62EAECC1E3EE7936F49853290BE20F9CD09FF0EF1638B6C8E31A1FF854C0A689F933EDAE0C024A364DB267B4C1DD37E2F1A69BE64EB93CBD2DDDEA56F31AC17B50A9CF9E96008E63583730453DB2779B9FFC4B906F2D4441924743B898F2C4EB074F085F91C2ACD13EBE8CA0FE546782EF36590C928FC1F5B2CBCCA1849DE4D1CED5FC27932565A9FAB5ED7D5C885A88B20EB7E7BD9E3027A8424F40A3DDFC4E1F0AB192A229FC56969D57DF61C0CD9F096B31473B8DEECB39D6127FABD604CA81891C825A192517152DF6BD0B09091D54F6314926F4DB49D5A974CB57B74D5BA2BE71632008CD7836CD312F220922E41D4A927202B514631B7A444DE7E2F66568B498BF1137BC988C72E08F1AD0FEA89F1A150DAE353EF2922BD0ECCD3A8F8E0B540169FC603D0235F0593AFC2E8B637A4D905E48D50A5E6EBD7829E0F90EA368CF1BCE340B1CF39623D4257951C5069943682764F447FA445D7364F32EEE39CA0DF5EDB72C0996498CE8920426833CE50C85CCF89CBC70678D398ACE430FF3102A82BE46D7518E32A374D00B31910ABB802B16F531A505F2F9BFE8E47251DC79FBA51F9ED8E832C25E829014867B4DB79FB77B9BEA8A1E63CFE1B8C6D0EFC68FD29C9DEC2F16B19F46B2D274F575A40846F12FA662EB1434195FABF19C51BB34C492E56360A3E7CD7EDC24921BFCB5D1D1E1F30072B884116AA225944CDF1332EA0FB333A7EBE61E52973E96C98B0E296BD5D0CBBD104BAECF0A1DA893871EB3E841EC867B8A8F70EC95502AC15804196B8C9915E5748D5421AE98DC5A3E36E5C1B06E16140416B39FE3DA9AC88C2D5D5B060B6183F4ADD6DE4D32E2FACA7BD3219810D8DCBEF4D796E9BB0E037BD22D6562D947FF9EEFEDD69EFF8DD38DEECF517AA2C880A3385851AD116EBBDB72F2DBDA8EF25C68507E9B315DF9A9298554BBA1758A56FE230B998A363955E9D012E04C68C7594312AD58A7D144F02F98BD0EDCBA5EC8160211CC609FDEDD425E494E4FEE561FFFB8C5D6AFDE4C04A16D93BAA8B89F2B159C1003FA0CAB9E69F20FBE2746A913CB0B8055420338A9EBE4EFB874D36D5EA0418A8C59812458E606B1A61E6FA6AE337D196944FBEC3DD6945D6459A8133557C1200C2DDD681A1761FDB9028C779E49CEC0D4E9842C36FEDACA5CAEB55E5A9E4C83C1FA7719C8422E2F7CF2B7D2D323B2B5ED3A1EEAD7632A62374B5EA796EB54EB4D4961D535DA9F0BB27DC13A97B560FC7C8BCBB7AEC2E2C7099E68AF4CDC25F1314FC98B34735052326A393174DF48B41AAE4EEE0768A2ACAE3C045374B7FF98A9336F0155B853DE1EA41479C148F32284A328F778E243F3EB8302876702A658BFBE28A39C428F540CF3C8D37151950BBD34A6188187BF3B2F494A8E168FFA718B8C1AB19CBECCC2E64AE70C321E67F26733747DBEEAEDB5FFCB32F2EF8A862B5923274584A6F75C38E11D8AB75FF5322E92C2CD2C267E3A897087037DE2DBFD8D0102FDDA902440710A7687CE05091AF5A180C1663C715C8A7212811C5A56BE8CEFDD8FB79D6ACBFB06DA4EBA7FF03517D25A6577F271C46D98ACBE4FBD30DEF52A8A82D63A1331491AB639A6806252D9D1138D5EDA376F67FCC9CA248C207480C6FEF02229FAE6BB4A0DA888721B632DDFAF582105C26EB2344979F41B85ACF10D13FCF9B33424175533BF04EB575BE526BDDE1CC3E9207EA16B6A8C1040304E0C4702B125AD3F1D5C670F052F256BFAEC836130550147ABAE85B324CEBA89564F29307EAC642F71171FDF638BBA5A32B13D05F81B1825A4857E9847A6E765E05F8B2190C8D78E63D2D5D8EFE25B54709AC60889A131E768C19A2C343C9129DC5F4E42845A48D22B2131A5DF9ECDB34E94DA200D929E284A038209B5794CB2CCEE4B2E05954A55FEDF1653A734B0971100E4A2491A0A776440E1E44E38156312CD8237CB3EC88E8EE259E72180B39D43E3156079FF31B368417950228608E88AB4DE2CE7324C400316FDFEE2983A47EB0F61CD09407F2559679C40627B8E907F958057D26929309E7C7982AE191F677D0A3A079C8E7421BD17BD0A03D1BC48F07B0A28C4BE1E8FA1C91172AFB89CA743CB3CE16259F8633F621C2EFF6853C381CB1A2D831B17A13897000BE41498AD50A8180A1DC066AB6538000BD8E9B2417F38287106389218D84E2AF824408BF604349115B89575158E81D93851C37217688C27BA5F06E68343E09D34B4EA3404BD5DB6C9E855EF393A5BCA80665BC0CC7856F14D500CE125CA34500FDE9EF19E7A0A319C591D022CD420C1656D09DD7525EB328FCDB0689A8946470180228600D5D0C3346B4637834685AFB0559CC07439E934EB56CE6B1592CFE4D57CEBB9024640901242B51C3DBB4BD0B05ABC6260C7D3D27D5EA057F215A5133F97989B2BADAB02957DD09AC700A1BD0C6FAAF60DA5031772B6F9AC155F83ABB3D926617750C54E42A0959EE3D73999A13978169F822C37185192BCCA836759691A465DA1D13C054C5E71E7F6C8F7A25F23409AB4CD093523E7F6D2195EF3782FFDA05069CF421F9FDC420D4D3A9923B4A097B6D643C034D4E4D46780F1CA166D9574EA63A95F5CB46AF77DF0626657DF2BA0D728FA562246B949AE1C89A9B08EDE2DF136CD193BCBF3D914F7FF5163C2E0D0926592AEACACEE96BD2D85CB7F563218C181E5669B493118FC3012840DE92ECA12E65E58599FF16A0030DDB61FFF06BC9D9F7112024EC67079595934F9A7D1C677F6AA66B9F145B1FFC70109246248EC8CE97A11E2567F5F5C55201F72CBE1F46ACB738B68517BBC930E0C85CA0E769DFD44FD01567850F742D2CD3A30135EB260103F889FE1B9B4D9A4EAD9C2301F1EAEB9E7881BC4C51FCBD39435AF6F0EEDA917FA6AD8E2DC8B2BCFF6903F34D60060078AB1617DFF24B39B67DCBC474359C9A26E382428F96B22B3D7FFAEB54ED526CEA1E0621FCBABC4B7A47D71E403CDD1BE030947EBE1A82B36ED8CCDF42EA0C2DC649120DE3A605B2930C98AC7966CD0D1D35EDBC9BAA91C8C5FFEE80C4D57C0FE44484C12D99E07490A639101139DF0B5BD8EC5A75C2F354371EB2D02C26128431C0C1C5450455D2FE72DE01F995A18A76BA105286030A00B6253ADC3909160EF4EE5FD5F8C63F454C783865BE30BE7385884E94A3A34DE8CBDE5A0A90F7836776F2C68A5ED45089FD519220520A454CA3A6E636CDBCF9879501189B8DE33D11E9CEEDA9BFAC2FC0F54A7D8412E81F58D24597C0DB93ECEDEF82680D82F4C2EDC4843623272DBE273D91943266617BF4F2344E9A9186AE71A5C856024568DFF250AC2BFD62C2BB2E8A88A371A2397C6199277A3BE22A5811896950808E02F064CFBEEC5FDC94397D05476280D6CB070E7E8CA7527A7EA1F276EEAB740AD7C94EF11D296F2FE93294BED03F207584EF447A5617E15EAFC2388954B9BA3AE9DC8FA18552FBCAAE3D7ADD7124D541EB6525C1511A28BF9A374C7D7F1E7A3B0ECDAC647F53F48B08DE1BF2BA3E722D2D43B0433A0658E3D8B4EAB77B7ABF3C2912B6E8A1344A5C8CA6074F369D761B36F2E892E57CCB094192DD8E23F05A09B0E998A3275D852058B49A6E3A6A8FFB8E9FFD9FE126170B12214A37BAAEC91AFD901D92F8E4BBB0F2F25D342559AF089483EE7CC92053BC17AE9EE73C39F211D4252DB3ED0655E0C926B07217C9554FA35DE492EFB79EFFF1A243A03910331BC267B54B88F6514458BFDC318D94ED2D1C673DA225F2AF8DB9449CCA4BF3410F3AE3CDAEB05B5BF6B26B705265E076C765896A6539B7984AE0DC1A1E686BB3D454EB9F04057F27A0FA9B82A88597ADE9692B04CBC67DC9900E819477D5921114C4AC5C8FAA2C9D3AEC64E12FAACCD9429F080CDC1B33F61FD7BB40B3149F71964C6E433EEC22DD8DFA8280079ACD2A8C15D1F1472571492C24CAB794673A0F5E2DC6340E2152CF4B442E5A101A2738CBDB655DB71D5370763069980FF59559E7949495EE21CD150FE639E5A1FE46441ABB64052443507AFBED13D4D90739B2467FC36CE0BA4598DB91A236A9A6ED4B8DC0738F6F294411A33E810BA6ECE2DE0147AABA32F73D705366F49C442A0C1CBE2FF19331879906DE55AE834E001F17F5214861A5C4891EB3252D159CFE4D1A40ABE2AFF41FE89207F6AD34EEC09D9BCEC94685572270B793013FC7D71346ACD2A9C54F09F66B3B7ED463B5A21F79C49121FA8E9D91216F5E86CC7B1BC754D8FFFD184CC83B7D18FAEC4B36365095B60372C5E4D4E80656FA965894295842F45C9473FA7BF3A88C8D38382A4DB1A0846A282D8CA904E83717BA8020D1C362227118891375B48793966B041AA0EB9D40E2E4A0133F00B69FA48657003923D071596C8C9F1A858061AC2E82A6D9561A01431E0B6C245EC82EE5D0819380B02B26DCCEE228A72AA067B47361DE51D6E61B3569F5B680F81F348F7FF047DD8143605D31E0BE1806779BA349D29C2F3BFBADBE4EB3EED053370D14A67E8F4B7C2006E564ACFA49B151AC26C6CC939CF6D28BEDEA33A3B84141DB41F532581B7A07CE05AF364BB7CFD65778C0D45564423D131F5C9AA1B13280C55D9EDA85081797DC57E8ED0F07617FC630E25BC2B74B8AFCEB937088A61623E5B9305902559A5899B0E7436A75A686BF7B18947041723A52B1C5023C382A9782F7BACFB717C1E5AA07540F448BD4E9ACDD95897F26971F13DB8DD32086AA6862A2FF8BEA37DF6C7049567EA61CB3D02FC05F5D211BF86C7E57AD50ED02C5E6EDAE7AF4514E4DF8FBC1BCA221BDFAEA7C2A3004FD338A9786F9E121AA400532D5CA1E5DC5B2D563999E4FCF1EAE2B0889B6AED5E34810BD5BC12841561A49E165E9032800BCD603089B99B4793E09535939444154CD27AF8C3236BCA12AEB9DF1B7F9AFEAF4DFF8D4CE51A8BBB6DF7E605613652F4881D5C23E515C77F80067A650089CEF9ED4B08BA15A508BC3AC28D8FFD661B96839EA460AC0CC596A2F5D586D1A78596AE232DEEA0D0BE3CEBA8D62CBC54617B7D4A124D938A2E5B949F244D818A21722BF6D20569FCE5C3D24FA57CE8CBA25BC100C35A679601738DF4C5BD2E5A6F08AC015184C82CCDE214AFBA2CE2194844BB1AD3519D748A1251BEFB4909BE0B5FC6054A587185FDDAC3ED8CBC208113B1AAF2B712A836ACCD0A81BC9470EEE1FF9F5DD655EDD61C57E91B2CA4F3CE1028436C051688746F367538BC53C4AD26880973CFA388F243B2A64792F8CF8749385332ACB0D40EA3D5C76FBE510E77C4A69C9E1103AF521F6772A5265F94A93C62FFB64C1EB589290829549576F819C93BC8BD7C74A89AD719AEFF6EC940073095186BA5001182E4F3DBD93E2FE8911A47F3BE1623348970A2F44D1C0D5D3AF1947B550F2CFF20FBBBFDB9B56D8FE0EE29487EB46DF7E6B47130EDAA9D77237562DC12730F4E47DBD296FA2A07BB333BF7633D753A6437147EEFA22E7FAEAFDEE813A7A28C94B86284A8FA32EA30A27EA7951DD34B88A1BD03060B312A61763DA44BC6588655D206BFA777529391F25D18152DCD73B88E766E3729E4560FDC51D607BCB6C417E3837D2C72805BB9C4A1AFC61DB437172BC9B19862DAC0BA377125F6741823247CE7647233F8B23FEE96BBFF450AD3D45C44DCA21864024AC77A4F7E7FE32CB5761B612FF97C18F63CBF39320DEB77690DD2E2C2AC64ECE6810B72EC676AEA1D9C3404102273B884413B38D4E7AF4518D64463C1DC3E9A23CABFE027ACB420066EFD4B7B6A38762CCAD1CC4277A300E540FAE1F72EBD556FE2C8E9EA89A4732728DF01DCE6DCB0ACCADDF807436B4EACED64372B0DB45AD4D298878E0081A180FFDA504CE01935C9F83B1F3FA820B26F15DEB8B391C883E756C29DFFDC99933A169352C3CD0E4518DDAAA51A11CA780724BE5397211C515DE240DA624ED80F96E8288C86BC2D1A08F66E8D108EBFB5E9BD32E8609E48980D4E934EC042D3433995374F0F45A5AB9E3E24B2C3684F48D09B4431F24B2083C4F26CE0A6493197C9B849913CAF8489CCFD1589625106A71B0D56FA49347F0F9207A2BF8FB7D10E8953D4A5A6A5BB29BA5C484A9BB9E8A20D216315E0CC2626210DC32D7992DCB618556033F57DD025C448D6E19E46E8F1C5604B2D0DC18A8549DEAA2461E9D5D3C2DF809CC571BA6BEA7E8FB5000FFE7F4FC53C4AC8B8DCDBD47ECADC84A06424C065776CD73ADA928DCC7BDDED721F58CBBDB6A1291B10409703706B2C85C4CAF81617A144BF12262CFDED33C203D749B20BCA3B5439CFE03746CA0E5AE2E5CD880829633C361F476B1BCF39EA1AFB1BBD26EB4F2B59C6F078A448CCFE3224F16F833172F12601574BCDC6F953DB6D1A60B51D83FE0BB3B2CFE97F397F64E938A2CCF031677CBDA8A1D31A9279A3D7515419762E1AD4F743A97501722991AEBAF04F8B4DD71ED1091B106320B0DB05C798C96B2333CE52B969DAEE0F8753663A41D7C470DE2C63A18A7838784D273C90479983ECF9A29030A71CB9B6D8231CA1AE4EF6108EF0E5510C710E5CEB62870281D8B83DE332B71E5E361B4C68F90CD66E03A2000B90644533F24DEB561282C06EF710E657788B3647E966DB7DEAF64679E7EF5CAEFF9577AE5AD935443511CFA39DB09DA716BF113BD02171E46E82CD9F29A96BD5CD97349255B2E85D8D7EA27F9D9A254CA684EAC5C97FE73D34005483CCA8C553EA72AA5982DA7ECC5F7E7E2E176502D87C26EE124139C6E37C3B8891890166D8117AF79EAA952DD0820075777FCE6EFEC78BB2413837C41C2DCA96569151048034381E037A47068C6D47AAA657184A2A3CB93E0E19846A7DB90E6329C11338404016397D4CFFB2CDB27EF63F0136760BA5751045F773A3A192DA88F33A59DC52E8491F0C39AA125BEAAE5D679BBC0C892643AB802067C008514E5CBA332E943FB314AAD21E78302445570D94359DF04C90CF67D16AD504392B7A12EC1A9754A9A33BC437E1E20BB5D8EA7BAF62458949CBC26C4CAFF7D978D920BD867F500EEF8548CD5E3E0D28957587F844DCC69D244F8366BA76F6A72A0824B53105E28540C024A65F500B7507D6417A7355CD8B030C31F2F357759F015FE71B7F25E3A6E0C76C8F222171E6FCD6C878B84FBD55F9E08788A5EEFF2BC901862384D99DEADED042F2E8C091A0CD133CF5BF699EAED41B98934F7B7CA74B0C86F68A0A165E2EB1558B5A687E41480B0461FF8230EEC6ACD14D154BE93E4AFBC829E79D9F3B7883F4571AF6C74FF4A08E9FF66DACB3ECB6B7F5FA9D635EFEF475665FB39F2E30931E8CDCBFAFA0A5117EB8A75D6FB1CAFBC2E62032CF848A59B6E01E498ADE6CA02130A0AF44C50756BA1BA0DB31D3E89A98E1E5108CCD9BEF26F1AADEBACA246CDC99EDD0D64E94157B0008967AE186817008BE70714911ED203998CB44369905DF93C3D94F583FC962C493748BF0B8F8F010DA5A5785DC20D50972DC5348CB42CD1AC12D4862315F52E40258A2D931DAA83B8E7A349AEC9980D0960D0818E791A8EFF867B13114A82CFE2898DAA2A7C521654570718D025F32297DE85207B60DA92610823DEB4F57D3787AB8F975B0A463A84895A3B9D726E59683DA731DDC1EB06416B32C4542FDCC644F68282D99CBD447131DF948C5791C8ECFE6DDDE1E57DEBB7F7406BBC1C53D05A4702BD7AE40D9F4513708EAAA734C2044F86D462B38C4E046A73A8B736A9115D966301A1EBE78EB0F8FF5E4B62F5BEDED97249141A4BFDE0A7039682B3AEECBF0B42191C59A441283C348B666E77E15131BDB87DBF1F844D6EE8ECAE38B236C372D786E4CC9422D17FBF58B5243909D4263A444C9047D6EC1B4C0DE5571DDFA3BDADE8340500B11523DD2589CFC27A3DF98F9E5F5F0D4685A0711B3798FC2AE5DC0B3FB967D487A645287A117B0A0F23A89E301E3454D8D362109FFD810DAE4C88CF87BCD61286D75A4E9A4289CA4E6086633BBF73B77FDA22777D7119CDB261C9F2EE7662824F00E8D0C3215BA180BA68EDB8A5C6D6E7BC8D266F02CCD56726B8F31A3BC350457DF170B33FD77EF2EB69F1D67D89F4D02F8510D860567B67AF2CEB10964865A9F7FD3A6F5C7B4901448F051F00D8ADDD31E64529E738B22844BD987DFED46AC8CF5ABAC6E06E91E39734322F890FD3FC37C352F500D83B5950A39A9CCAD1E10618260DD6DC66BDBE6B7F6627D11E4C0BCFC4BC240E9EBEA6D4EE4DBCE51493E88722E0EF10299D4903148F90A1E2422BA95DAC54F261ECECCFE94CE0ABC6D46D21C874D8F56317891B66BC31F07E5FA527D02B5949E7839C00809941D846B93D3F3329CD87582B8925B831177C021D95FBB02FA3B8F58BA7D670990305767FED54BE6ABF71A2ECCEB6701BC31FE8E3036B0FA87CC608D98A9624DFEC71F3E988165BFCB013F284BFAA16C44CE846B207CF484DFED26E1B8B59B1F7DD69ECCA5D9238054E2EC7FA034823033827D3B544712D36E16413F012A39EF3DC6B5BE85221A659150BC337981C00091F7D1E537FB51D14B1EF9AA02DF917F1806B4A35CB7F57F601A7AA902978CFDC755699EBBE54ED292256FBDF22001FF03266E2E6EE7AA5FCA348CDC09F00332B4FCE6C369DE6EAE36560541B7EBF580925D3D92E7D46B0410D3502043EF17097623BC3A83DA54446BF03A87E632EFD36B6B4205C4C32E10464D1A49F6EAEACFBB8E1741C55532B228E3A7803D94B85FC601781C73D1EBED743171884301B279698D3ACEBC5F4251FD8A2424772A723BEDE482C372C4C0CF4A11130AD2A3008AA805B3B3BA5CA2B0C6ED4CC4011AD45995031BD8DCB5D6903BFA11C8E55595AA062D2F5263BDD8B550E0A691CCE327488864214E66C9F2232A399FCAF35742B55AD3F25D180E090C47768D834A7206690B24776136F3DB8AE6078ECC909770C99F0BECA764B03CB6CB76EFF3DAB417A170AA909DF23A1C10DE08F08BDF2B306C3027A271E174E3CABACD041559EE4F1F05B0B87631DDA1674FDC228C70554B40ADA103B94450BCEA7C3B11606AEF69726CA8CF58746E4CB558C8A850A207F575CF3602AE507AF7AF146F72DE2E6E31B1B1AE5211F9D17D0DBA3659FE9C33D98E47A30AED18F9C5BD93AC741F77F20D0BDAD23B57A3A78045F1686520658B099640213B037FF66E8623459A512CD1BCD9A62789EDE1B4871EF875D32297806E9F1371028EC83B5FD71FDE9329A2C9BE9789F39DD1C4F17EF19FB3B4F66C465D7E3A2C5031BC750C40FE896D4E6DF0F783E8155B2A9DEBA13949E4F07AA362B26DA1DE2076A515312771D3F33D65288832AB003E131460377347D461E055958BCB0BE268D3998683906913C128FC2A2E4281F8C8B4C3FC4609D3D016506C598997480DA953CD10E560BD3A0DBB223E7482988AC63820F21813BCBE6051B6BE04EFE695F6618FA2F4AF74CAD0A4D83D7902096350A1FFD9E2CF0393054D8009B9979A6B3470FCFC3DA69F401745CD29BFF3F13FD895DF38743558894A630FAFCEB54842208B4F7A9915D855CE6C595BD8681E7D22EE379FF569008A1990479444F75EF15BE183080A503DC0EE85C7AF55F40A6DFC7CEFC5BF0BCD2E3A0B6DBDE4ABD9B90E9FBBA952BABC0B792AF820BBF7563C92DC16BF9899619E8DD01FE7DAA898129ED5227393E1CD34CFD2DF430251D5DFBF847D565505CD4E97E22737C924C4235EC6CAEE7378BC62A533EBB274ED545EB56DCDBBB58C033778ED22AE5A2F607E7BE052022BE1CE43FE7F4DD4620360950A93F149A9802E148E389BD076987630A4D94A39D74EC60507AED911DBE34A852B76DFDF98DE821CD915C4AABF521CDB4ABCD6814FD848A1CEFBE8DCAFE8201EEB78D15CBCD51EBFA717D67468649E496E70E35F0F899D6F8D8690E338A7ABF9A9DD851F4909CE169BF8102238C19164EF5EAB2FBE735BF93242D35E0B027542079AD21C3FEE57D980391C2A07CA531DF94B94AA0F22A4A4D0E3A1AC31BD34013ED1AA8CDC72A48D1756A67E093CC461198260DEB431A047F5545C8E83761AB2C0EB92F15D859FE3E8162D615BFFDD4F85FFF8A59D6F52006285D66FC6ED8ADE4FB9E02025C7F6403C7862E2AF01456A830EA220276CA171F01C7AB3328701DBBC094A366B660A6D7A3BE0F1B8EBD899DA47D96AF3DD115438429531209049FB06D3DC95A728A38B3F3DF4C40C43486E8F33D691ACD8217CE218B51FCE23BE018B31670DBD6E3953FA37B1E719539ECD4D999912EF8C23E31AEB5B88FBD091DDCF2C696DB9F83ACB584C05BC016096E42C9B2E6C32373B1E49089EFFADC03275DBFA2D58F8B17C40A0A1108FE2DE4246A3CC7B176D0FEAE612ABD6A9F04F8D07FFFD09391A4AF5C6030D948A963ACDCB62189628ABB6DF75AC4F33519A78EBE4F284958947979B896A36B0E2DBB76AB35DFC8108C0B6777BFABB7328C0AAD592AAD6FA2E04DC76BADC62B6E85D2D5379AF9D96D0578DC95B4BC47B10F4EAAB2CCE5D4C42A68D9B8A441F1534E271DBB7CFED513ED2B9C77BC2EB0E0AB2A025D78ECBC79FCAB905BC456E9531C57FFD9435AF245D6CB0383CFA53ED685CA3A524B9297549F4FE982F62B1B8833C15D59CF3F29C19DE6681B34A9AF5403C79032A5F00851789E9BD0E0CA36EECD32C589BE506DE3993DE4132840C41E2ED148F257D5843F881A5D0257C2E77F802C721AF7D300C38D9EB17C03EB2AE7935F689A5ADC1A940F8395D112D4A988125FA3B598DD427401D4F6F4C0A08214779780A51F6F0B652B5EAF4E74B7E5E048FD23FC44360FAE18CBE66E3748F6C4742D4F7AC0AA294091CF5F54190AE5C2E8D3CFE1A042A29146A05B9158E408629395C8FC8A5633B01B56340FC2E972722B02CBA8E87E6BB91876563851B3C03DE2E9B94F603ED1DA45D7B25D7F0C47795AAFF7704B1A28AE5ABC0DA192D0CC2E4D3399B7B6D6C5416BA48E1BB5EE9A261E64A980C0A7B0BAD4162579479579D369E4B2672F36D45F312D5E566B80AB76BF97F287FFE08361660AF1B0C18D97B64A4E07F659BC52C0FDAFF52F87704A843EEFC4294791D179622012BD82AC413AB9CF8BAECA5F4CB934EEEB82A506B60E7F201B5C1C5BF11BFE3DD88B5D58C9CC1D1B4513C0913CA624949E59CA7CC3747A72838CA88490E53DC431C896AAD2F73B411C650E0B78FC2EC89C99DEE380D7BF8212364F9FF423C93F22DC477CDC3D3C0A25453A9657748E4E7FB25647BD58B69959943615E9A0561A05CCF15288B2030FC1506E9880B6714BA5CF2A79A9F2B3A32A03F774163F58F8B15431E6B8739516A51BBFC148C5141858DE0FC397B700F775BDD25A7FC6229814ED6C4B074B620CCAC4DA4FE7839066CE5897639B72DC633152BEAFA850B01810A509F44746AD4D085610540C95A23704BB640B48D749509F7FC7E347DFAD7CF8304F4508A539B9BCF08F968FAE9A74F8DFB4E99B233E8B60621DE8168986CA66024E1463A318491F0C5E51801C8FE1555D9B01D8A2BDB3335386CA08EE0EA9E7918B94B7F6F28664DDA1882FDB288A52BAF2C2E97A110325B81B647AA9926911480F72550D35C9DF969489C3CD2B0118044C994DCB1025029A2CC0CCED0A533B774F5B3738F005F0BFF717086AD8C12E905339A7FE7BD29207558E8B2157549BB2D5AFC04643043846131264B89F81A865C80404B861632CEEA005BF1E0F9414845692EF979B458A969F8808788172798A6EC69EE3D9AA4982E2543CEB491255F6D5CD9B5530E4DC8B962F6341A7C75A21BA735AA887150B47455D624DE6BFD448F57DB9C5F0564D0FDD076CE96BD7BF50A090E81FD86EE96E2B5117B753ACE0BB53EE55F952648D997F4E4C3993C15D8C2C0E967517CD56C7181B2171514A3B9717B1665E1C50C5E4C3ED97860E4CDF4EBAB74935A276CB57400F4610949910DC008A7724BF31656145B8C2558EA8C32796FA597A34E0EA946C0FC0F07D5FF79DD5F545989CAEABFE65E1615F48E2F5C0558E90983CAEC33F1F8D03E1BED5A3E5023C1C3B1B1669944F041F343EEC2B3D372C18065DB37264C65B6F92A7743AA02CAA3B2234AE6F7EF7C70F2D75B52C810345086D94BC89DDB339D174FD4BC106D661A478745652A1D12022FAD07D30B3FF5B573910F005AC222FBD604FC24AE571AD8FE3F12082A718B7569ECDA375559F15B9686555D932717F977CF455F0CBB97ED7ECA7A60A248EB5B742DAF8CB180A71781ED2E532017ACA6178DA60400EDC9A7C34987755A91B5EB238E1A19F9B11B1D1B83E6063A7856AD6A0BCF268B28640910374534E260ABA6550F41245A9B33CF189A9557C65D3C5DAB6E21BE476230D02F0A347F1CFD8E28215E3C40DB4CD28383B4EC8DE7AD8044068194ECC4B7C8C01B654A4404BC5F4DD1099CEDAC809A3AB3D51FF5BF5466BF7CEAF08655C3F60C6EB60FE1F1A18CE3B7459D732D9AB005FA80F57FE28B24FFAF4B674D1A32D9F62FF353B4DC3A9A39222DA84AF31F99E94684924D72233B245B83563C12A394425AA575CD2C2834B23617B5D710EE8FA22B76EC482C59D252C06A288DF81F665B6857468B5A714FAB7E96EE0662A8CFEFCF2C82D7154F0C75DD6E5E9CE3144D887DE2B3BB8C5B4982D878310E8AC504DF7FD3F5DBEF66D4855936DE35BFB8D516221F9E22A4A31A304B0EF052F99A4AD0BE61DF4A5C5D248F75AFDC0B392E4F1961947A545B8DA787C163C199DA39FF759EA5518E9B5F720ADDC99BC5AA489A701D79CD7B1C641B30CA34DFDAA85CB7C10D0D51894D08455C3B291D5ED34445AD47475CB8EA85CBD0DD1CD2E4C626CFAD92132874C2985EEB44BB3CE8C0C39ED865819409816173919DEB9EAC00A60EA2C0187C05314ACD1174F38DFD692E2B4599415768667AE0DBE35E2671586688F9048D8D61C03198C8951C61C07FDACE9BB4130EB45F344F8A31BEB6801F898045D69EC57472DB814F42C55E77D39D2262BC26841F0262F373D0DD3807802F9BED7FE5F27E6A7A50C44ABCC73BFBD733BB6FF5079DB59DA26A1290539F1EFD2557E24D33AFEAC0EE1D263B16634B5A66CB55F7C1C248EAFB861ED9365F059F781E2DA33D2E3AAFFBAB05A3C6875443890B7AFAF68BBB15BD194F5512300CF10E1EA404EDFEC4B3A6021D70DD3A55ED799C7E84296619A1640A4D0234D091EBCCD78408147A3DF6E876736BFD8EEBB1ECD38FE3A5C27EBAB4A54255A46D1DE621EBC067EAB17EE0A57B1D4CA61A75A315BFB966063E813BF19C184E833CE265B212335CD72CE3EC23F1DF6CA026EDE1D441ED303C537791800B7F04B88D3F59FC6FBDE81B4C9D19275DA3EE7D646F1DACA22FB0DECBEE3E00626321E0B1B1D60190212EE75414B8A4E3C04AC87A8750497CE876033C902C812B8C432305590247967470380881EE1639BF2812281D173A5653B6E2980FC613F479B4A841EBCE4411BF383DC435DCFCB23B16F5357EE431095B8DC0C2C6AF7E1773A3BBC8BC699456F712A48DCFCF4D6368E3D1D7CC3A6874063B2F9C9F96F6E5FF5F6AFEE209DDE8841B675FECF4E7D215A8A22E1275C4BA3693B68493859AAE488293783BD6D3C61E905E04E5A50E0738D7751B97FEE76342A7F9FB73A2B96CDBD0DBE541C4873E54C859B8DB59D1DA9805C0E849415D17140F1C0ADA0C68F438C7741639C697885F0A7A4F9EA2CA90E8E63B213F6537A45687C1F7E8EB8F58D225D19F51EE1C020F7C0ECD120889EC3BFE2C746FD721078AF262F114E253A235FACC401FBD5FF0D4FECCDC882CB7A6093B7D3EFBA2DFA380710680102DA0CA57BD31734ED6F8C29DBC57BA582335907FE46121FABAED4C0E8A213C46ADAE574024307BB04ED67F99413DFB0E29C080F4EAE72B284979E9BDF84764CA9DCD71E88CADE804D0A792F618E5582921B3B0C9586ADFA99F916D89A60FCF6CC36247F1EC80D222359CD63097AD9615BCA0675840E57A4D09E92CDFB7BE54104BE1F0B70F599DCF3A75107740839F9080E8AC6C47F6E5EBF681004BDBA3ECAC2789D54BF1B7AC32671AFAAB33D130895C4FE7A6610B5B62E454D243CD31C959AA4ED19402BDDB70833A920D0F52126E1092389638518DC1C4C7C0DF58C3CF55F7E11930AC8B4F5A28FD84D926C2DE4AB06E2F68C027B285F4BCD0474EE7E7A6C5501772ECA9DA5E34E1DAA7B4039BBC6729D13183E055B5E2E42E09A4DCD04676165AF9102B2CE27EAFE958B42A4DA64D84DB7D4A922BED536D9FF583D91EC6197A773FC5D962B13E0388681293639B31469504DC6DD4F5DC83CAAC0D9A86F35DBB0A2AD6104A6D8185E791689C5CC6DC286024EA1CABF30CA6589ACDA40BD09A5865B21EC1F3FC175BC58DB29E60DC8FE25C7EF64798DAE83CD6628472DC7EE73154F45168DA535E9363700D729777ACDB23CC3A422784736016A17DB9C71861FD206E718DA4CCCC5AC38FFFF0700FF374C79276C9165FB450FA8718A04987950600BD1941A873FDAE375EB07F6AF67731EDCB008EBA9135A9C7EE795A4294B8282BCFE1BCBF105905BEE7143DFC94FB91D53A8E1DA651803E115183BB5595861FBE1D172DBE97ECA8C47E4CB69CE43E5528DF6DEEAC30D2B90AB070FA6273BC30E991AA46F99C1F93FE3CBE2AD5FE175EE2F953838129FD427A48A87EF07CFFE6BCFCE8AC310D4B7207322B767B160AE6D1D26BCF29968717B6ACEE1562FEE3EBD1DB57F9BA4BDCEA99FBF42ECBF9446DD6B8900516FE6DAAEEE0605E9EE429BEBA62876E063E7ADE3FE04432AB72D69C48D47B2D86BBE5E424551EA68B9D2514D17DD76FB3C777589B471F669D1F15EABCEBF6B251D3976B287DE37E75351B3A482F607B4FB6E3749324DCC20CBB7CF4643617935181344D575551A4E4780C749A8ED91F64D44354C18EC84FF7E028F98796B8BB3F9BD1F87DC29C86F1659E6C33A639269173DB4AC23A1C3E96B15320FB220A288384D8C2FB2902F71C048BC7A0BA891883AE843934EBC9F0528BEBCDFE64589C1530DF762B53318EFA2D91777099EB68DA63B0C703473B440B01C6AA4BF78DE360EE2CF90F7638DFE76E2DBD30170BC8F21091264BFB5A83A9CDBA0438B6CF085866A443FA6EC15FC1FD7B07498CADA16330209A800BCE37381DBC9AE5CCB868DCC28D48794865A065C9D4634201C36058E2942740ACAFA84C36557B4758913FC3913B4A5C9FEFDD2E8031E57FA373EC79D8BEA35C44155A51C164BB6064B580F8105419E748FBDA922872E99C0EAC21F1E8CC6FC74217E276AD9E87B664845824B134408BAE18BC044BC64B2C1BBE1FE714F769AC2253141AA782F9CECAC909AF5D2F7EE195455E283B8629FD00D4920D0F59FE91EBFD223D1D945AB35CA7DC06221097A5259DBEB9CEAC09E59D2AE8A9346BA17DB038D8F69CD3CB7D1BFA50982E22D9224040C1AD4CCE2F8D1296E312D9C263D5A207C8DF039F2E7CEF187DD8E1E0EAE158114D1FF53180A3C171E5377879816B4AD4689C58F79D9401F73B3799C5CB92C7C27984703A59E4AFBE629F38FCE77C707CC2E63915542ADE4F0F89B829C6DA0F3CE89E34D71A0AA11199463F2214589B65AEECC1FC1D956F344F909BC0A80E08243F9BA48E00C0CE005C00A7641CF4DB4767AE2B9B6BC0AAA7DEB326F574CE4795AC0B500D2358D38A8E408DCDEE54E48CD33A44225BA0996A7326E4EED33D466EA224AC59F56DED57F8DFB52E3AB399E107A6EE2D219D54DC7A993D0F1EB57C3DF10C87147204F3B6466F09C41AE1A3E80C488CEB227C67E8531FB464DB9129192A7504C008215C925FB24878E3A79F1E56EA4084058D09353FE000B5AF8EE3DE0320A936E20A00D5CED5C73F123FD57BC88BFF7A42563F8449953D70A970BFAE752EC3EB21E856B9F4ED958E411CF06D0DA370EDDE77DB89D017A536735896EE2A47B7B95520AE44FAEC0C5A2E34D52EE9114D6FB31B8014CF8C9423F360A7AB3BC385DDDF54D731FE1CC6AF4AD89F823A69A622D8AE938250C49E10BE7C2AEB1E444274F20198DA2238A0EAA895C478DA0D3DB43581641C01D2C23F788CD59EE6B91D90ACAA2BA8C8269D95E63F1B17EF8B4AF19E8A520DF67217AC727DFB2522F7971DA582547BECA01AC2890F06E7E4C653B8D51C3201FDC7FBC9EBECFB93ABA6211B4665C9585E187C4011D5EEF4D74DF54A8C39932CE06EAC79496D7484D3916886B60C1524892B3B847AA7B690040F3EB87E4ED66800DD5C848C08422EB9007F2276DC68BB40FDC43F6E91C6EAA88414CA9A0B764B7ED252A7E756CEBBCC2ACB8B89CB9B5EB5F64CD7A263DC9ADA8E0510D6CEF90F8862CDDC1935F1CE4FC43910347DC7B1EB8C8D27A7E511EB2216793194F9D65DE95E1E6BEAEA5BA06220706E6F8BA95343ECCE8B8A5229E33DEDF51FD23CA8181675B4196D6639A94B1D8C2B4609E977E124C4B5153B4DAF505945DE9C40C86C70095C20672A93249F1A013889D1E391DB5491E3CD5AB704E5D4C009D65F385270AF11278A8E577D97BCB2FDFC51A061319348316790752D2B71D06F471105D2B45C1EADDBA1F8C9F7FFEEFC9F1979051D287552C2865815851E56D7F36DA8AF2F902A864ADB59C29480ACE84C3FD3216B136152498A9EC6B02B12D96A9A77AFEFBB192960ABA100BA4DD7925A3A706F9275B2AA81A0632A126B2131B73ABF6652B6FD9027C1C02DA3F379A3914C031EF31CF57899DB85DC7425A3C5C51071D87FA8B01579D6E779B4259A44AE656C7C839A69F8C83E0907DB426414BFFFD8806464BBFA074307BBE67AFEFC382C8C39FF341FDFB6C851CD2CF4BC1A9F4EE867740A22A3CCD60C296BD72D2EDDF058648B3ADBD93E2CDDE1735122055D687A390A4CF9C73FF9221AD3532C4C2212ECDDC79F723490A2CF27EC8B589732D9E2B6C4BF589E5AC430A8AC376E03304DADB763A1CFC3B57FE59EFC799713C4521324596D2B24374631F5E82BC0876C1358DCBB40C72255AFA60E60AB0FF37A32906BBE9E0404054544FE31D8D426BE6FD8CC1CF4E67152C2F714B11289063BEB6EE1BFC69142F1DFE1FBFAEAA872C941A6249F7090A45D1CC30571FDD35D32AA573BDB11471874911479D1EA1E0C18833CA4B7387B4404B5EF66B3CAE57AD323FCEEA0FD302A370966741F255D750F52274CCF8A170689D8A5CA51FB67FA9D5CCEB065E4F4C93E72C509710DBEA1DD45B6B79D24DD0CD1F0922C9F95C1F57F320F510764212066CA92810BF3A2C2C5BDC33BE374792146CCE67AEE1FD16F703818C1DEE1CFF34D4A1A16131DD1E8330C5AFBD5F5DA501B7DEB1DB0788F7AFFD5348B3815623B0140B56B0126924A17CE2A726DBDDC89767E5D38A11F2DCAA83764670BE7B9BC26AAB33906E99D64E6498766E0098E5B6E1719A9C7F6BA15E8C2173389D93ACFECAC2584CEAB24F24090E336A2C1127A50DAE64BBCA8E63D0FD157A4DF9A5EC567A93017BF00695E9DA97789ECEB408F9A47F81CAE671E8A601283297353859479598A173CA6C9A98EE8E735484F6484658161A771CFF625B15CF5BDC1BFF99E08CF7F8827E86079AAA77216576608720E35C91AFFAAE3FB7E53AB81B82F84A2D7A8C2E74FBD1AB0A15612DBB20C4F9D5A52BA1A82D5BB220BE849D75EDE154A778EDA20FB347513ED3B60F9DEA2B3F85FC38384B58540D9DD2FAF6EDE8B6B439FBCDD32CF0DB86E9F933A83C3A4E00E3C74D404C9F93F29F5DD74549664FF3C453AFAB81F759DD9CBA02AE0E7AAA31EAF578A7248EF3D349763FD38FDD752027826C350991C65D825E7FDFB992FCD8ABB8157300A606467FA309C42D35DD7CFCEDAB182EC85E6D0B2764DEF8314F8E528AC3EADE8E352AE8E708CF45BBAF3E05821FE381A3147925E03E19AD5FA21D9C9E7F8A83C85D4C16C368ED34DEB67355C2E8940397A85394C5E45E3EF79D9B79546406A62CCCD49BD828BDCCB6A89854F0E87775F56D69DFA1644171A2FE966C668B60264D783E5F6FA3FC14879F1F4107BFC946730B61D01CF13B86261B1A2BB3330554E166BA688CA83EA64AED646076F7DF9AE4E65B3F51E084462DF59F231A0ABD8923549EB5B59436A3435A0957BE532BA004F30828AF2023F3EC92BA1CE9D16F22AA00B70C39C80AAA3616A4260DD31BEA9264EAB354390E614966974F0B4D6B666CDE25B940920512B7A93DDF1B9BF156F86781744707E655B129FBB526D1CF642DEDB6AAD036A23825F8910A4528AFE0659664CEC2275325E77E7F82FDB90BB8D1A61F2E875EE7C6A71656FB624E5534E1448141CBB351E450AE5BC516F649092C67FB3F28207C21B73DCAB56D8524C52211646B862986F886C9D0C75BC941A5F31A8F8FBC68E9DEF286028BE1634D930A9A9333BE2FF92A70A3CF0BBECB19C0C58E0FD8F6E55546EA3AF70AC372BD37E7FF5EEC33A50B5C74FFD76D548AF5D751EA4C5B57BE15B42706447EC6394936A90AE8BDDFB8C10CBCEDDA87F609B577C1C642DCE6D4E1149B976046BC475C3B7F15412FE50C8D24B5A78318E80D34A61C8293A981F1D70E9826792802770B45A14F36750506F2CF1D6D0452C56B555D034108BD465C6CC1DA0160C1E8D7E18E6013CF71187CA1001DFBF265E5460746F81BBA1EDA67528D8B8277118D2F9F163E75AC9D959FE955E1F3FF336B7AAAE41AE5731DEE9367DD793D183EDAFD99618B95C680F143A4A7BE7A4F35BB1B968E496F8B7EE7DFEACE4F7D48E30F4066E4D6781FAEBA0C65D11AD72793C0610EE47EB2BAAA3398C7497A266521074E6280BA66C715815E6903F235FDB579641028B71567C1F954C74BA372E751B08C81582E740C468D69DB20B1CDE01EC64F3717D393192790DBE4F0DA56E68F41D7C6725273EE21C7FD409D003656F960D818E883224E1CA0AD315C73133E6D87D4C014BA04E9493DFD501FF486E785C4D5A6C20B30F176D5D29D602A4369F8E5268E5C5AD179D94E3FCC042B1D15FC8915516D4D0A999DA6CFF1959D3D1B03985D31CEB92EF6CAB166639CE25FFED072B6C1020586DFB508F4CEFA2A01D005CD11204A3038D5DCCDA6D3BD824962F360CE7E9DA640AE734163DD7EB4D026547C37676486FF76BB89E53B4DAC2CEA4B4338E89F48BE877DD0060A05FB69BAB82A695923CA6FA8F93717759A4B7D4F499699F7922D9BCD50B18C3E9DFAFF03D03AB22664C0AF78A524542D685F40CA1DCAD3583C5AFEC27DEB4ACB49C8A2710DCF8A01180534DE0FB3B0CAE23446B0D8D6B3995F14CC3819816CA2A60E888C64E4CAEECFC0D668C186A20779DD6860AE9341E333ECE17D5BFB7B3F30BB5A0693FA84DBCD575B8DBE8C58D05F9A3DBE958E1A3ACA588517DCA36F80DF728F5CA6E98674C07711DC0931C12F86DD9626AFD7C22B63B922F0E248661A70A60FD02BC5282B694AD39C3CDBCDAB352C9399B83531B06C84A0F5E6A01B690B0B1564B1930488AE97D3B1CAC7C3FADCC96083BF4182EACECDD5AB4B567892DF8796189CEA16B2B4B38D5FE9C4463DCD088889B055A3CD3144903A454DA0CECFB69BF5AC16DA365E95910DCE1112365F49F4B2F252E18B6A80475374D758EC4768DDAF405D0CE4C1E9C75C1C0068FA426E162996392283BDA3BBAF561DE75668F789B6BA2C62DCCFD1162D6E6D9E38B23343B4EB3F1D302A8B9DD9EB775CA2027EDDFE4F1B746AA14FD22FA2500309BD78296B8B7A6386256FB84F883B4892F9625DB2A521DBB10BD7A35F65EADC578697F15E14385E5DDCC8EE1BDDFF06DB728E18A3873FFAB5D4587B4C34FC5B89C600C8181B9C823F169624ABCF29ECD3033EBF1076A48952675407B922104CD4636C2DD53217C8240EA999DCA86DCF025510CFB558CCE4423F48EE47270C27049AC65EFF6871F6F034B439009C86BFE5473EE826B1B1074D4AF5122884BCADD0A43309B45ECFBD3DFE0BFEAE116C767C09A8AE465BCAB8ECA63F915DBC5591B763DF8651C8A7B1D042744A1A0DDD306F2F394463396456D57554F3BAF6CB2F4D722D76CB22EA3CA170AE47E7209E33AE5048007F0B7D03EDA3D433326AD591E6A68972FCF8F3797EF8CB08ED575DD7DC12E6F94900CE3F98B9CCB0A83A5077556503AA4F76E23762202F4F77449670BFB37F78D9EC3512F54F0CA98378410B9C225E24E7AF2A8F04DFED51D667918848A17841C52B2BC2EFF63CCEC608E02A097463A45CC61F5FE607E85A2B35BB2334061D8B8EB47D3E5D71943D402D0E1BCCBE47A0649FD118FC523B13E17EC4DFBB0A99078D552C67C27E18C4162C4A85C4B2AF04C1BC925014843712F671B1DAC95BEBED385ECBB5114D1C287D4DBAB97C8B26B097D5B5A95F117B1694668A366E1500280606495D35540BDF49DD84C37F9F01E535EB8FF6E3F0D3236E4F65162348F9C862298C01BA81751C53A787762985014CA8CCE8EF88AF864F6F2684970E7F7252F981479A415EA48FCB4361C52C5289E7EE49FE7B5E76AEAA031FD7FC4FC280E74E32C2E655AC5F532474AB3488A4040E4F33022AECD13535808339E5C16EC471B1357B65A48D752A59E88F5947F5F1022696E85986B1AFAE71756A3EC03C6055E869E1BEDC66AE4991F6DF477986F62E210795A3AACB8908EAED3F5E06E4376463B0D6490CA8860011FE92709CFEB5CA8D9ADBABC952F255968B71E994C995B1F47049C128FD0C9C588220D96CE36418A546F2DFFDF568FF4EEE72D3C48EDF77E975F9794F5DEA289A92AD5F76462E196422B54BF90BEBA4D1A116F1F1702B9DF52DBB7C90D4007D5E35DBB860F6A6B52E47CDDAF64037102D8EEA3F5AE1AE42BE91D59703BDEC67F22F35A1873F1313CBEBF3990F99DB126BC15D347E1D2C580F7F9DE3DBB1F031AC2385002AFDF00710AB7BBC221ED794B36C0087FFEABF6FEFC38D57D020C0D2B5347A73B1BFA8B6E912A9EBB475AD8FF0C49DFD5872D3414C8971354D0BC7EBF24756C9ACFED12A576FBEDC1C63914F53894654D712FF03276805D4919808AFE3AE9CF5A9B742812E9C3AD0E02E94ADCABA22622C91EDAC36EDA5BA6EA213BCD715F870AA98E340C129545D0EF4438C84EE12E901B8423B4F06CAA829A2F143594699E2E8708922769CD85459AAA674BD224A017FEC42A6AFCCD32E1EA2DB5CB9F310619CF1E95C06E8FF2C0EACDC74B1FE54DFCB7BD3B7399D561EC65C8C7BE88EA323ED1E68F2C4B078D851A91BF91ECBF5767A12D152C01EDC43F94C5EE2AC8769E8438604720BC918CAECB779EDFEEBA19D77A75267BD4572F16BBACAE45A3E8F1FFF423F3D1C879E46CC8337FA33C59D74ED05BFEF83E5CDA1AC9FDBB9DE8E3B089E1CC27BC415406DAC7811116557CF428FD0406E203C8D4D95E00F812EBDF5ED80115E5228699B0F6759953DFD7E6CFD1159CCB47C774293CB7474DD800BE8C91A5CD7B630053232D87A438288044CF64B6F7774D6D4DFC63908F4328720E57BC850E768298A3F0EB6E940781EEDC98A0AE5AC84A29916A93A34629766644667A0EDA15FE73E11CDD26C6B35011DAFB9F2E25FA5527B9A6FC0D0C5F35DA042AE208BD5ED7B71720F846CA2F68C4DB6C5F457C596F8A9A72D1753CE5E0AF1C8D51C84E210CA49C23AC85AF82D4C27FCA9B768C1C06B3490C4546D58F1AB1EF1727F8B6757C580DEE59D4F60F7BBC32A595396EDCDE49BBAB1BE9A77DA0DD9978D4FC49B18BD2F881C0E27B8A22783EEB4E041D61FDC8F15411A742F197AF6F81570CD032F0E8177E34CAE9DB07EA4C4E01B26FDB2786F0551DBA4954265348E1EDBFAB3E9B3535289970D1A67706E10FF9CEBA033AA286E0B79B707D09B67514AED057FEC807B924821078487F24B5B8057A334F48BD2B0E11778981515C1027574E448A38BAF5CD516146B9894198606ABAD74DF92B9598E09E1600F95D546E44384B26CA4FBEE54D01794B69CE404491016BC01AEB080A9B848EB800FC2F43F6BA9632435DB7964C28713523E5CC924721E3D00981513481E698AB47FF796A65221A007ECD4167BA882F2B048A41B9CFB9A3DACFE5A8697515110A59907792CE805791E3518597CA9ACB2EE3A3E62A6F1A67A1CA850FB91C3BD1DAE20E496714B40063F1EE40EE45EBE4351DC3FBFF0B88A1510C22759F9E43070DD1097E1E88FE31FEF19A2735779EA810AD6870168FADBCE8F330544BD84D55540AD27C8AD76D79F5D74248A40F6F29D60EA75D453148BEA09F33931C3F9CAE2DDFD4AB2A0F653281106D2C130D69154F22409C9E84A6CE37E63FDCE2BDE5E15483C4704CCCE5B230DDFCF844220DF046760D5B69FAB84A1CD13ACA4C2CB50A70DD82464544CD0A1D135F156EF03F613EF277B6B8EE428F919AA1E0CF712BC819AC376CA8F04F4C011AE25F1159D446E522C310F2BED45EBAFB7F44CA99FC975E9A5D665C569EA3EB412AF28402615869F9934A227A639E88912733FE5CBCE14F4E4EBE7671AE78244C9ADF03FABC3A52E07B81A995E59C2B9CEE4A9437A52447D2B827C0ED0819369206319CC9BC3BC82D83F305E07BC25EE2FC62F260E866C756065ECFF33A4431EB770B80C4FE32A7E62836060B2D0364B862FC09B98FC98F5D4E5DCB94CB0A6CBAD3D8DA09390C8CA3709DC5AFC86B3741AA276EE69BAC8FD22FB7BD4395E750AD08724E9C792BC49F033144017852A670FC5C1BAB9F10D0222FEDB3ADE3C89382F327F1EE4B2E9BB0F374EA843115A682129EB22C6E5C8DC73B10EA53DE665A4564004A88D30B771FEDF7F1F1D82D9426DD5D5D12D0AFE258D53BA0660A1518AA8791DD4F1CDEC958A24FDDB36B98F6B13B0A91038961685449524FE9D889B1F525DBEAA225AA779E5F087F579E7BBBD641FE062754D1D573BCD646367BFBAB46275B980CBD6A4EB6E8F57365753F5DAEBA4EBBE46878775DE43596D3664C8F7AB541F07504FD7F22A49A3EE3011F3B29B79F85E2BC5B86780872FB8FAE42E572E98481404BCD1A1608E2F5635F0BBCF55F9BB2DF1E7F04EFA486480A656A2ED862ECA1198FB2E8B0BEBE2E8657EACE2E058462E705BA802B25C38BF7D8F00695A545550922D3FD097F6F11C26D094B40FC8BAD6035E63C14272AF7F046E0E32A357041A9168B93395FDAC93C7D1BF4BA2F0DDBE29FCD71532CCAD147E7B166644608664D2EE62C54B1BFE334E9DA3816AFEF02CE268C926CA2A57026642D572FDF3003D5AF7D3517E3E806D0B38955485FCA6E4364F1B9D787291117D7BD4AE24CA12DF7DD6D0F8C7F9E6E6477195FBA43F9FF0943FBD77007B027A843769DE975D15A5EF8E2F3352A88A15E23AA034394894BD88B4B2F3EC9C4600BEF1BA60FA58C5B71BD18ADB9D4314EF6C19B0CD157B9AC1E772BD70DF88469D1F05CF7813B3B6B9B4C63413427A09F89FA199BE8B968874E9122003A0F3F6563063AD9CAD1D6505F4C2AE8359C495542222DA9BEDDB7B8C93C4C6AD4B334C71EB9048E509FF3D77D2A949EC94A9E4A89163160D51890CCC00C85CD917ABBEE01D5F394618FA812686900BBB05AF5F54837D740759299FCB812BC314182DD8B0CA023C70A6223A8048CE9A3B41ED5A28E56C8E2F942C20F62DB12A11CA9FF0BD764E868D3A68AB261969A1E86FA568A2C053363DEE4159C8234B277F7C3F8ACA356AC0A8E71E3BC2C8951BB02076F0CE4D8B92F008F4C76A981272FF4C6ADAD509F0587635DAC7D7EA168828C3471C0EE6A7B884D3A0C95DA70AD768975CE8D680F76CBC912FE27B55D0EEDEC29E64A850C8CE832D080E2FAD673832F7B9E77D380DABDC37329AE77CBEEE33E2F6C43F29E64882FB0CB783A91DBA34A7B4DF4DE38F0DD10EA0526BDE0B8E0D7BFEB87C2690096F825D0CF4F798E67DC840E67269789665E176C5DA2BAA79F652F971DFF74A6144AB2BE96B00AF12760CCB91282D9A36651224373D814C219C83908121C987155F81B1BF0BF8D9504BEDB9A816148F259CAC86AEBF4B9A51FC1405E5C941B0C20C023A90B370CA93F6449F62D4B2D9DF77D5681F704E31E70004911CA3A71CAFBCEBFEEEF921AFF30AB5B249DA765BB6DC7CCADC782E2E1CBAC31C2AA58850282DB1E58674A2B682426E32BAB7201F66F8F4CDEB6D0D0F5D2EA7C5AFCCD841AA2646216892B81E207A8B0A3C1762BB52B8D8CC94A0410985747091852C919DEA9374B02B6EFD7675CD2C4AA2452EE4F81AAEA65CD1AA0B5EB54F95DD26A563DEE748CD545373D0A2928A140353E043A9E4C67DB48AFF7A9538615E68801D762DD08C651649FE3FF6737A217D5748C1C65D8AB51A6D8EE1363568603FAB52ECDD7D5C84D612DD4C203984C0564F0D0AFAC3D8C20026D19AC5E5B824460B23D93F1EB423CA8826B9FADCCE2E2EE4283E3ED2B1B0747B8DC0D1F620E2F91AFBAA88706B3E4702DA8F8EDE61D850913D544E7F2BCBEFA7115EB5C8831CFAB31F7850FD1DA0CD76FEE77E3DEE4B9FA37E68C46F1EBF0B3C963DFBC5BA4F359D253011FB2E72C165233B55123C187DD0A1CC1EF0E17D3552DB6BB95BEDBDF1DEC8B991C95B74C23F7DC310B2809980EFDAF37D1FF69679D9F1D071C7D5F8B4EBC0DE8E3C7548E8AF20C1E9585E82D3D9ED624B80753D79D5C891F2B84DA1F65370FE3951B23799B2517FB3AD7BF7E95B2DF00CDB7038BCE21FD833B9F1C1F460C77A8A913314A551273BBA40F69B6C8D1370E6E32BB6E0010C1F8522CA17FA267AA8563E4E18394792F40318A7CDC2774B13BD16253BF3BA8BF4144839D06197AD8B826A87FA0B93EC68A5767CD249B27AD5FB51C2E1B670B1D8695EFEAE794D6455C4EC88C37162D9475E7036D52457F2F3491552E90FB33C12F7CD1516830F74A8CF35093B9350F8D1F7C65E5C3A6F94397E30CD8ABC4A4BBC86A9C011EAD8C25374834C546A398194A2ECAE9F7740A765679597BFA7024DD4540E5B293382C4A44F33EF9E9050684C50A74AA3113F579863237C1F4C221621C1AAF6182832A5F701CC939677507028272F869567894C608BD9524C1641BAB195034AF5E95B1B22709F969314AB2B5E76AAF4A0B3DDFC9BE419BA623E373908BAF81A3BFD54D1B526FA5B8735B118426B449A5DDFC086E58E9F5870D8B9BA387E226F4119C2B1A74BF97139D36B174AC2DB79D9BDA1B35121ADA5D87306D84DC8FD2628AF95FF37200A7CFF4B03004A71A5F5DF5C2690E9D7265B4B23C217BF12EB8CF9501254ACEBD9AFB241EA51DBC21D41F4F77986D0680098BFE06EC5DAEE1388C2706FE232DB5C6EDAA01DAB2DB2F5C14B5D6728CC7287C07136A739BCFEE2FAD82E168521BE45714ABDC8323B84C924CC61DF006E11690CD5719DC404B8193A096E2A0A1A8A16729DC93B40453285702D07E835A42339303D4C39CA3E2F3FAB8DF60FD58311683D7F746736051E9BB16E53FBF3C17E4ECCCD8FE3B5BFC844A24261AF5D438CC361F58FBFBA87F4E90279DAEB05CF5D4581E5BB6F2AA6D5EE8E46CB2C3B2FB8F99E8DFA393DAA022E592FB3F44B9C01E07FB978E3746AC63B7C719F8177FA9B517C52B6FA2637F757176BBFC4842ED828A5B59B31269E248D4B5F75B58A330D5B68C5213AEA7D6F343AFE140F8C7AEA7FD03DA0E5059D7CEE0FD3660D406631669A8FDA502FE681400FA6D7ED6A89D690AB45648C553332CD89CCD2078744C257EF32A3BBE767A09E2A94D3EB52F4A8FC7AD83A6E74CF38EDB435D5BB6B0A1D23109618BB1521BCB871872C2121C1EF8AF58DD37CA512BD34B4D58A8C8E63F3E68B0AA664B9EA6974DDE08E9D9076C5B2306F8676DFC75450F10A362F42593AC62F61AA69FB03693033DC09AF7036CDA436125B149ED19997298AF77280837F54E0FAA4F351C6BE478965F5AE55C9767853F0AB44DA3367C28562FF76B043D749E0780DFFE74F6133467424B4818A4C09EC71DA15DDDEDD89EABEDD115D9E324BD333D794252214D6163395DD43E6CE04FD49CD204B2839831FA3D3F2C0A59395EB78620184C8CCDB4B99CD5B43F6D9EC9F972ECE7D873AA62DD33D3559254BACDA190C320798210EFA5F851CCBC448736C5E7AD0A48B4087755038C64EA767F751C58FB24DA96DCC488D0736C8AE8A4BBF2396C1D33F33B3685D43F5F57F3EDBDD9EB355330566D7A0B597040B1F8BDB9454429B3FE31230FD1FF250E21369C194F121A4CBD1559BA6E461DE412F09FEF5CFAB46EF87AF3865D5D76F16BE2C56E6446C6DE7C9E2DF23F1DBA7F827204828C6FCF3A1223F243B385A7F3A3EB0B1AADF6958C4BACA6E781AC1CC1E876455C3EB13EB657CF978E5C80F8316FD06E6EAD50987397584303BA9B7B8F487E7EAF09C1E1F05E0447ED5E2A9AB217F6B9D81963B774D1280D9A2566502B78F8B6642E3D30646D60278082D7C34B9DD6868D2157BBD40401C1545FD710602D570C82C1CDFA101CC3562B557C1328329C23876BA9BD2A59D30A438EB52045CED72A09F2CAD3B8934A48C4A49D8B3F2F84519974B2EC5A3B4F8C9ECB29D53251AA95B144B8AB3628E9054606E22D1CBFC28A7CDA44174E4984C19D81602CC0719CFBEBE4FF9288F983BF0FF174818ACB1CC22CC76F4A1A9AC759C3E3AF56B62FC8C99C9C4A604136234D6AA5FA0B17AFDA216485FCB32CCEAD7E1AA1F29262E70D277C0CDE82F8126031443824F9544BEA43E248E64C03597A2F09D18810CC71093F67243DE10DB77C1E03336363024C3B8FBA2C135D314BFAAAA674FD877A4E41E6A6ED1E0C5262BBE7E5615A59064CEAFF862133206D4A87E7A908910CF956F35ECCC88114FE5F50ABE224737B73C0E93082160776B2BF66B2B2A4780AE99CA7E101AFB871211ACE4A6F170C285B9C16E8A43F241E2661A8ED2DFCE8AA03BE5516900596731E17CA5BD0B4A5C0910D07873732B967D0CA126BF39F6C73CE1D56EE9252233364A2981A603613E8656A3B1BC3F817D177860CB8E67DE33E5A66D07DFC3D3F5B255A3D9169E8A51B0964240D2F7D9EAB8D6B2301984100E35105DFFC3AFA372AD9ACF965A5C382418A5147DEF2133887A1DE7B7A655707E8157C9EEA1D5C7CDC5E1D4ACF852820F403B654A3073A115D51016C6A825D436C3394A2B7F43E0868C9B9C34C670E588882854822282615E286AAA5E1B665A62F76AFD319BCC27D49F332155F7B4A91AE4DBD7B1CF33BA74887A0DE66ACABAFFFF68D568F9A199FC39123974673C131D427C5735E0D622E7115FA0BB23B811376C809C607B7AA69F69F869C44406FA4346A6B239C95CD4418C4ED7F860979EB6C1F8A4AD3E9D744D4C0DCE8C7593259980B654A0DE36D092C7E4B868FE8B67B51CE5204A429AAB5FD14B52D517CF1EB1F74E4A56B846CBF6B0A6032C9FEBFCF728320B685CA121EBF98A857CA262BA604EF8CB5D22E2F51C76D8191ECB58B6B4B905BBDFA398A2674B0C7F5FB9E53BB4647787B23053CDC66AED653237D0E98FFD6ECC2107D6B2C9920E865E97EAD832514FB9B5D387C271ED28F59562BF2403B9D56574B2BB2397E9E69B092DD154471693BA986F089F05C438A2A54E29B432F15AE472B05AACD4F00EF992AE8821F0CB6910DDBFD4B2B3925C3E69B035B8D12A4A35122DDCF536227B09F1EF33660026402A6E7FB5FB06ADD2A4E1B55C53F64766F7C8931676F8132F3BB38C5E406AC847991CBB8F4EDB988E2F7D181B5AA3CC19AF68B32631611A5A2DDB2109781EDF7230B3FD2AB614373848F489DEED96E937854B4D7211954D68E2BE42D8978282E31051C5A03EA5341D988B0D478BD4DCAFDDD18090402839D23BFC6CBAD7485EEAC73893C5C87F28D96097709C7620446023B9722753327FC9505B2D3F7152ACBA405A6C738A8D38FE23322CDDFCF8B9402C3846E912A50DB88F0755985538601418B10A35C9AAD3D6A85FCCC61675013DC810115EA4712A7E6CE7B7EF054A14A65CEB3BCBECB5C1234D6B8EEC3E9BF52C7AB93E031275EEFC0FD40333FE0199275CB39E9919DF683D377C2B77B9215152C2EE7721C26B6B5459EEF4BB108ED9F293F6DBB953644198861D80F3FDE36C9269A18CE04F71B93E11D35AC015B6E594D4AB496FD678CA5B69A140DFA47AAA4EFABCF66071E87CCE268CEDD8D1AAB68D0F6A026557E9893785733DC00916CEACA14B0036069F93DDEE917DBFC265379D1A948C44C97610B28A8F6658C3596615F23BAB6F5A7082F0966851F5874F858AF215A612E6F8AEF06BE93344C9C9EF8C1A69060A3392275D4029EFA81951E27EF0CF59D68DC5FBA80EFF70FC7F6ADF1061A02CD48CF01F612E4143BD5554C313CFF09FB9139ADA6DBFFF15B8B94D638CAC8B288C5CCF2B9364ACB1DB856F8F685DC4E41142D36159529FE7E14460BE3C6452F41E427834FE4512E958488056B0FF5BC662F4F32CD6C05302F92C31848287C60442FFED397E2E425D1703CCA94B38353B3C56E3CDF99D4B09A6F2BC8B99F0E9B3511CE7482D2AC6DC1C89DA66F11B85A4847BE9CE96CD2A7F75B7C8A22D891C80EEF2A2AAF95409326FB35F69C453B71BE38C010C5390E0BAF7E4530A807ECCB2E637A3E8234DD0048234E60130548848AB0D593989BAD1C93A7098D6D63A7D2832E613CA357D2D197039C8BD5D2BB8ACA8A38688BE1856843B045385F1AA630B519AC145DC404BC554DC812D9BA311188841CF5FF37D9E89F0491334B784FAC4EAB18A4298B9FF9C8E9451D8E76EFBE5E7180CB937BFB89BEE339E1FF2337DD777F0D0D7645BE9AB762B57B92A059B181F225C705FED12FA1C8FD5A9C67F69B62D1BC7F9EB423C9822523C0BC007E84548EE187D86AF94D77D7A0E39FE3E9C2D084A49D0787D83085C554317012F93234E4F6E3570F193562C298BC74B0FDBEFF2693CBA14DB233347A44EB7CE18E07B20C94AFAC0550B03FD288D434A8305106E6536819672F1BA674EBFE9211C12AA2C7BEC8E685A67FC7DE8B51824287929685D117A907DE3B3E5058D553CB9CFEAB7F3C009A5BF727D7CF45DEE16D94FE8A91D54A13E4B6DE9FB20835E6FFD15760087E81B36804DA1D1C1CB7560FE18C8075AE84B1E94EEAEF4BCE2F6BFE7DBC0F3F46BB26434661F3372FA6D36A791798974FDAFEDF929FBEB9C61ED39AD17D41A41BCF38ED9A6AD1EE6543E17BF02349FC4DB1DD5B134526E8E2C24B661964ACE16FE856959A2D8872CE4FB7E40CD143526AB0841EB179AE2F6AD3FC485D4EE0D6C557D4629C053D54E854E014263CD67AB2BAE9BCEFDC2F228909AE29D1C19603D13128CDDCD5E7FF0A21BBB960CCF39B46C36B9C2179116204FF2682538FB63A17B67497E75F50313E274C677742ED3325347BDB693ED5A56BCBDEA7C62BFB0BE7D3FDDA536259201D0A06AB5860276FF2607DCC59D7C4C8D08E921BCF0765EB0A71113A7F30021A5AE9AE365B7D19CF52AF56842A92FCC9730EB48252E77D22450C09E034EE702EF7D1DD16FFE7FCA201002CB02CB5BC7FD85BFDD6CEC582014791B504E0ECC765BC8B0C35C6CBF35C0C5B61ECC0057B26AEA140D81AF03959A45D8205853F67A99477BF98C34F5626CFD17ACC43884508BA22C9E313DCD427DF99957AEAC6ED308694163A772EC8193BFB7B8E3D47BD3A3CC8CC224DE37DC89D90DA5DAF0A2B4148CE60E4939E295901222202D759E25986F7612216A265BD00D28B3D9FDA34379003E73201EFDA6D859C0DAB432F275ECEFAC642F5AEA3E27C1E204E58D47F51EA3D3928965E99FFE3C483A499C37C32B5C3D5164438CA299C182D837DEB92F6E534951593D679094F1F48A08F43A5A490F95809232934D96394F082C6FD96E7D566594883637852FAC33A699AEAB5A7E4FD572588E7DD735103A43109743F4BD0E76326C1DC0E2ABF041C0C00E85463EA0BB19A72C1BD42DAB9F5F293AFFE0E166F5B8CF8ABE5FA7A485AF6C4B0C3344FA48F383C09FA46933AF7B797A37E55A0609B8BE4F2875F3FD5A4D4925076283CA9C285389A95F0F8628FDD691D80EAF44C6E2A5D554BD3DA50975C086198AA6378B64F8ABE87DD65BBA8D671F2AD579A99E2034238F2A1C6C7D443DA7D0B8EEDEBD3382D1A4A9FDC99A3EFF4B8E4BC5E166D15F428DDEE4D0CD2D4A0AE12673153B7D2CDF473A742B5405ED264BE0DE404707838A185E29A4E6C70AFFE5F89906E2DBD2329EB7B4168B9A8C9596EE2D338028AF8490200CF8F02C26CA15D6F0D0DAEF77422923E06B3C3BAD821088EDE48FD388DF9E5CF7748BAAEF7FFBEA9C23BA056D6AED16920A392ABB3DE6DE85ED77BC53A4C395713A3CF2C4C43A1DD11C9F9E764B98FB53A9E37ED0D1BE9F4F3CE76FC8929F42E5314B5DF8E9C8B56266312D4FDA5479F4916271AE3A04B85424373B119704A8A9896B8894EF1D5EE463F9F6ECACEF8ECA1458D8CFBCA2F79AFA31B17C89FA6E687F2E6C0937ECE41F4168462D38AD22B483E59884C73AD6264CFAE427265EFC63EBF05CB47D4B19D0243E10D49AE7CCD2872CCCBD0F24F957DCB4A10A753F7D815170813BC044E802649D8E0C776D75F4D78F3AD6D74145A3CA383BE27DD508F5005E0AC5DDD2B77CFEA5F66B535C1B5854182C05079FCDF454418C41D9BF59EB424FA78563121140B84F0F5CF106F0C08011FA8E21B70CE5F071F7EC49A2CA00409C39C80A97A2D20426FC2A44FB5424BB0B703D0418436B057DA0E4787F4944E437253CC682903C152B353B15DCBEBA9C623A8815BEF8972A716583B4658CC6876703CDEB00E9F0BDB80ECF1441710C2C319BA42CBE631104E5ECA2A235722A85AE69CA5CD5AACF1B537E840F215E1F1A58258279FA1BFEBC2BF90634C45FF1B1F8D2DCE7598957C23B2B50F6F6E8B300BD9C334910635357A96F4C546D660F4D600152B3F966F6E548F64C03BBDFC5413DC15CA8CF7BCC96758B33EFDF86039705549772846E9705E1F2B83A0E717F84F5D0EF9E8CB33DC294CE39C469CBFADF99EA51786DC923AE2E75ABEB934E05D6F90670C67C2B4CB456BD8BF0E5CC6285286B23A1D0243F4012CD99428A83770F8C6DAAC7C0ED49FD4D609910FAF2E2C99E8C084F85C24551840C241F670FBF8E93CEAF036549F8BBEE4C2CE6F32579E7637BB9A55AB0E47460CF9FF4986704773E39995591081ED79027A185EF068ECF068C0006761EB7CECA2866DC7C80392DC28F542C4094263C0013E4DF806B81A7E22386C82CD3E853615EAC2BD3EF5CECDAD60F146B25ADD2ACF5A50C6A22BEE0D7FEADBAB6C987941A80B50E9B7A6DF4BB3C9B2D1B36DA0809CF31AA943DB9E158CBB1CE14B6B89040439FBBBC1B4D15773E5DD87BEDD4012F088816EEDBCD71311D1FC9E29E4047F1809E6F5B5BAD36DC29738F0CDC8DE26313EEA5F1C40E0C8965CD1015A7CBA35229D9706745ED82EFD3306B5B48C50D81E796A4A582634E428521DE564D4D4E85AC035B1662D7351A3B89F532D6355BF25389218E1F141D6236C8C9446A73325D85C1190A9725C8A2480E6CE8CDE741BF26C59673B6004185A007642C75F3A33AC38BE112F4426AEE179AA831EBA76D36DDFA0C75A66C18DBDBCD675DA50399A22482F31845031B6D003CBD1FC0265A491B8121AC8953D05F2C1915270D2004BC1153EA0BFA7A5234281A9406FFDE5D8D104A661E01EC2756AEF9AA2926EE62E34EB778CEAD1F90D3589E24C313E772CA4C46B246B2C07094433EDF38CBDFDDB954538B7B36B74B6FCA01263FB01D62DA07BA247D061D591038717780867CA13703955EB7CC3890161BB7BA2236BC0EDBF6785210843E8645EA5FE402B1B4321858B587174D4E131772D993AD5206A53BB951F7CD08C458219EC708B1C73B0A0EEB1AD758AF121904AA30D5EA611CF063E72C28F463A63E64B91895810F59A2A20B2B2F3A8EC9ECA2CE6C5C07B71BC32DE8A74C2B33F16DD6E65784A4759C320DECB128795D2E1DF6EDD7A7790563ECB47F6DB7EC0A96EB1687B69412430A05498B457F0F205372F020C87D49EC3AE11CB254A7C2B838D503E24A2814DD352E28349BFBE480EE75EC7695A5A15012998590BA7142525E2BBFD3440BB67D46396A55AF677187C2FBABDCCB0755C81F03C822413AA17931446857B7F40E3C94C458DE743B2CF5768F8BF983D31B9C7A9EF48C3C5F7AA2B4C6B83E26FED4EB8ED3423D3158453EDE29DDAB03C3BBD4516C1ADF673564CE89FDB3D14C88B0C7399F619A56A266BCD904B068968402D715C8F1439F1074279C0D4AC54691D5D450CA3381C54530E7F3D3BD0D00BF69076F83F6528F020A2C76221056AA24379A435DCF2B435CF0F61D07A42E5A58F81F338962C403992A5DD81CAC6605224628F7A7782E497892591BFB49AA694CFE7C23F8E091BCD91A3FDDA06ABBD49600465B829E5DF6C3A082249428437C289C25974A3C26BE027BB66273BBBCD76A7484F51612EC159A1F3D44305DC5B4897981740889CBAF4D328B505085110DADDF095E9B5EF172E1B1B553F2C6596B59E1F6EDAE54A83092852438BF925A75267D59F90BC0DB6D32A215097AB02BCA756B960F169E660A4FCCCFB20E91F0244FEA82CA63F2F701C3253A07CA00D2A0F3778427D3D6FDF71E0D92CF0D26DA087C9309A2B78B9D49271516B53DEAF36B4A66FD9C6CFA31D93984443663AD358003865EE9A1E6E4625F9A0A1A793B7951D43E14657A67CA7177CE8C53258C6779351B73C0853375E0791F008BDCF300F2028113A114A956118C94CB18C512F2B16A8449E54490C5BD6811F8EDD1C9BC21928A934DA68D851DBBE3D6862BF69F6EA6EF7C713CAD4DA6C4900867EAF72407C3AC2C76643288D64D781E50079842F2E751AE6FC7127C28EE9FB288108876E7F0A5F40B69833BAB630E176F211AF702648673D1631D56715ABD4BD18FF763F5F40079072641F5416994E1860527745EF6FB4FD3033E3FE9F08CED736D221EB79BC4BF40AAFD988ED8C0DCEB5E8B3D359A39624D80244DF708B8C13B8718B987F525A2B21487FB50CF041D9D199BCEE9175E4117E88B178948DDEF2E696A724E2EC78E41D3ADDF0BD6810DEC7553DBB137DFBA7EBB1054D92D8F667C91D58358EBC7BED4539797B1F8EF28D18BA229ACD82E1EE6B79CF531562796C174BDBC4F0C54A8ED50B63DAD5A49C5580F10392D2948543A86E03E5DC33CCEAC033BC2DB4843802056234D5DB250DBA71C01A390DEBF215389C3E092F67C1203EB10787382F2E9F4AE534E0F740D13C7B2C898B4001C4E32544AEF40415F4780D6F69400E866FD47C6EB49851354EF1BA5C2793743D6EAD6FD804BF12D0E05BAEC8544435E0C5D0FDA7F2B6CAB2C01670418C7D47A332F747EE5B1AE13532AB2B49BDE53B358B54418084450C435DDEC464C933ECAAD61105B195FECC59A40AFD9FE8C31D5760EF26758C75276294B2774EF2124D2BC2C17535D78FDC43C2C8D59EDE1E939B356E704D45FC655143C86CBE8ED0A19F078FA184A9154D0CD45E2CE3DAE4A37F36D554819A3AB88D9ABF30BF312AFD73550832B2A722F958AE629482DA1BC538E0230E7114E26B268A6A2A15769AB60EBB84B6F80BAA82CBFFED08DFC747F19668F01860D65B0DAD8ED23E60A5A207EBC753B67023BCDFB64137B6C3FDCB73420D0694CAA0406301DFE54BDF0EEDAB50A9D673120BD92053B54804B54287F7D5A865E094EC52D5331E7F71D7BF56DF452C5C9EF95F88376A853BA59DEF879EBAC883009F425339EFCC84693DA7FBC0D915D9E1C146130A8549FA8661DA6F3A57A8FFA3714F0F4143B0308A8F3C2EBD6C89BD78EB6857F63FDE89E0CEE04849A43501376FACB93E8'
			},
		]
	},
	SiggenGroupItem{
		tgid:               5
		testtype:           'AFT'
		parameterset:       'SLH-DSA-SHA2-256f'
		deterministic:      true
		signatureinterface: 'external'
		prehash:            'pure'
		tests:              [
			SiggenCaseItem{
				tcid:      39
				deferred:  false
				sk:        '6088D71F743AF2D1080A9991C746F46FB5E5D70B41D5081574FD3F302995073F3E5589053D578CFCA5BED79843A13346D15D891EC1A38FC14382BE86DF3626F2373D4566F9E290681BC84535EB2E689548EA49F602060271B12E06A1E44F757F213666ABA6724D7AE8C18B65341707655CE4241C4AE314D798B7CBFBF7C0CA1E'
				pk:        '373D4566F9E290681BC84535EB2E689548EA49F602060271B12E06A1E44F757F213666ABA6724D7AE8C18B65341707655CE4241C4AE314D798B7CBFBF7C0CA1E'
				message:   '02C25B2AB3C9227148AA5D1F124C0A1D318AEE3016E3F257EA364D4B9C421E2D017B0456A01B8310C49E7839360E3A3E155E0DF355E1BB0618FB4637DAE610C0E4942E4C8B1F7C3E7E4412D2EA0A52306D2831AD0303C22FC88F751C590155D6706244893FA767470C10F6181083968E17A0392FBC8123281E6DF4F267884F755C225581996AD1A758EE2E272BE09CBC82DDA4A977B2F9C6E4DDF4104FBF363A3722F8AD40196BBC49B0E2B5480706127D43B29DC3879855D0969A04271A573AA4772F32F31A00357B67300F07C95D7EE21B2BA6FADAB26755EBC8414EE62479C0E97EA586E92EA9EAAC7775EEED4198D7E8EB4B941824231CB51B21C3EBE1F3DD1EFD48613466CE67BFBF1EFDCE1C700D8B2C2FDA0197BD32E0DAECB79568A9CA75440A5D4E240418C54C2CD65603F7A2D2B62C95AC6821285B9786397E93B4EB957400C6BE43C3B8C1DB4222C018C966136B4B49543F3F760AC9A011DCC5F3086FEDEE1F6A0A0D1DFF80D4EBDE2BF1FCA862FE729C23D884946AD0CC61C23895C7204EB21472C912DEE76C2CC3D3E0DB9501D4145BBB29BE9F0391331DEB056CAD97BFBF0686FE7D775A2EC5E17888269EEEB7662FE52D87E0543912EF406C0CAC4EA54BFA7FC94C6803FA89430912D91681738AF8B1BB52E3B93ECFD3668171E371CEF4519EA71278AF18EA3711411F240D7970B2507E7B43'
				context:   '19A520D0F629545634F7EF551E8EAAEBD3117468446057BE273AA2CFBEC5E0BA6D21B77A2E56F69DDCA0526BE28A856960E522CB761B74D01F4F26EDC730F78662D2E0A4F80AD0F6DCEB83B831770D4E2769FFB54B428D4DC5B085FF4CD2885F5983E3F0D8ADD3609A6E0E03683981A54E72BF4F90500A46C3B852CC6A6B64EBEEECF1B31D5CC0E7B98F0555885005177DF06BB0BE774C4A37004D99948DEF9FC397546E51FE95B9237EC7DC9B41461052E75A5A0B2782435B43B2B316E465816CA097CF6058FED74B76D840BBA78EE9B3637DFA0E5C405B67B5C650D6E130FBBF8284292AFA74D0E168B74B82EAF82193889446DF2403F0CAC2CAD528E040'
				hashalg:   'none'
				signature: '7A0749A428A7DD2FCFC0A824D33A5A2E157EF49556E19698FC310E51C731BBF4FFB615270640162CB645655C5338C1F901CC034B825ACA79F695F87725760AD94B7DF19800D7DD5382D0E9E80281947F2FF550E89762712F59A6E33CFF7261122368DA17379B54AFECE97DADB1C7526FB626AFEC24B349FE0021C1B18C2EC6981F80C7F64D4FE30D63044C8029EEA061B80BABD4D7A752119AB5BABBE1483ECAC02E36D6BE248008EC2250C470A11427685F34DCEBB730C6DADBE6E45EDABDC3B94F8B8BC55B3854CC0D1EA5D78A0884198BAC06569FA461DBBD05E520CA8EC6DCA44FE1EB917615174CB1151A24EAF13FB0F6AA3D592DC3D91426F704D40C6164C593DD5F4BD35CDFFAA977BFCB6ACBE2CF10B544DE22F4E6FFAE7F5CA89E94429CB0398E48719B22291BCB0EF8B67CB845069F4B6778916B869CDB37C86BB586D5B4F556A4EBA27CF722C8538BC1B291A9FBFAF57A0C39902CD56833874F2A572CA5E6A2C35C2E2CE5019D18FA4ED5BADEDCBD8535722B9DB7A287C09360ECEA4B332CE3AD2B1C2A15BBBE34BC5AF132D2E5C6219394FC3E3C13A53265833C961BBA0CAFAAF1849D1AFD80597CB799802AF89BA5531B47DFA5BD85B0EC3FA1262E3631CFF1C03A9E03A33886113502085135D4E8B025C187381420749F5B9DCB0921C0168D25B403D61EEE422725CE5F23360BD028D93EB3BAE72169D1371A24E6B41E68343375F0B60DC7D0D2CD84EAA00E45BC94EFE8D5886E6048821FD38FBB024466936EE1761554F3B6E69B874F85E47AADB5B270DCAD52B9C6B1E2E935ED7F21A14106AA57EF017D8F170C7DAC684651DAC32F1A37C018A54EFBAEE60221590A336E134FE9402FC13BD3C8369FD979A4B2971494D4673009F5837C91E56F3646C8997F9D9E7EF973A10C9F7C15AD7D51BE14DA02083C016EA2EF0367A7536AE21CC57F9D5B3F763D5E020CDEBEE5A04B2C4BB1051A217001C331B002D736F6D4BD0C4D2A3FB2940C7E344472E0F78A0DA73D833D57EFBA0DA2FF2D0B27687F2A7280446CF15CFFCD3D6C0D76F66BF0CB33EF7399BBC01D5CBD7DF0EDEB31BC7D35FD7E10D911431AC58EFF9BA934C532544D63F91ABF867D51A436E3D472B3897055B77A6630E3C618B8C0F9216B3359BE7CE1F7B72A76A44BD980DCCF15027DCCE711087CC3E27DD6CD48BFCA5AE9CCAAFD0E9CBC54AC5F4F3A9194286E81A117266D4DE7B7352299F972E5DD6D757DCCB2E096366595EF981C26C2B6B990F0AE1D5CCCB0D42731F913150FFF7F26BFFB98D37B55FEBD92BF062810CEADF5F44B68EE1620E8898CD379422B0CC8F72564146082D399511543FEC64C5C3BFF0B8169B2ED255E84615BB2963015A8C0A4FA82FBB3398769DD4C9F1E2A844AF7AC597EA92B9A52E893BD0EBFF0ACC616C50BD9F15E35AAF73B8C91985D1A622C32ADB045251F2D174D266785C2E1CB5CC3B09AE3ADD5C13F4E4BD153BAF87800EE724350B106451DCF5BA1EE2F1F4E58535408B86678C7C7D378984E87E4396D54C46D93E4FC45D28EBCFC7838F98A697AF3714AD81B73159621A28500317737C88D89F3170DE0B0383F8A1ADB3C6B2A83E049BFDFA39A48C9623455748253D51EC2B115D9D2881F60AD5D77FC95179F0E8203FD55B102FC233C8AE3D4B8F9B7C17CBF7B9599AB3F52168A1E5A11C158E95ADE2FE4F30A3F8777286548C16D8A3D41CC60BF0F38719E628D4EECF895817B549160B9F4BD848B53D2C1E77D98235914AEDAD174BBAA3A13B2C96A230A01FBB5E7B6B5B670EF885C7920261C9CC732FA2B272E9841CC96E2AEC36C08256DBDBF15CE25FCFB5708C5852A062A92309B95D171DF40E9FABD4FDC373C9732B211E64D7C80305D5140061032C843CDEF79E56F418337AAF24387631EEE4D182115D647B56AAEBD94A7537030B1D07E3D6BD0FCDA146F9A7D2E86EA4E13161AE858D884A207CE2CF4D06ACDDBA2A144C4D22623C36D7331FD28DFEC95C51F7FA1BEF609B7EDB0824BA1A9828CF1B586C5F3E1200A3DCCFBDE85EF621ADFA1445BCA66AEB389CD8DC8D44CE4EED836001DEECEAE94A633A88615AE0A3C5E09ECBD6E653354EC2C8713ACC6DC38F124A46D6BE0A8FCEC4709D8605A63A544281CDE4AC6B45EAF8B5DCC808DB527051F81A1A69B0F57D70574BAA68DDCDFA74547E8E5599D90D8B7D6CB05B81DCF223D502639C3507A52A4551A41317E1A871C6F735019633976DEE407A5ACC50DD8C415664B5AF17BB91D684B23AB284A31A3DF0C769662F47014EE3893946E38E711B0DD1FD958F08BD525BC84DFD2062D4310EE73F7F39799CBC096AADAD1688C4125B574149601E6ABBBC47880AB2105C137B6B73D077077F9269758FA36EE2167AA7623FAEAEB54C7E6382987940AF734966F69A2CB9E75666CC4B2A6BC641450DC57BCFBAA197AE890ABA3FF1AE5B356A410DDFD56B0899B139F00154A5E0C6D8BEA4B902F2421E1CEADD31BE5B4632A84C46FC06E883E8D5C3A5E956E74FFFFD3F9EEA14199A92C70C8B12C505B80C72B6140E3C6377E6E4CFCB1EF5E86CDB86140E45E8C14784C179B8E2D3ED79FA4EBDACCF4F4915815C624BFF1FD4A6B334D717943B81F5A4593676600CD8A1E73DCDC1E41BB85155121CA52A1E5CCDFBCFA87BE7268ABED027086E89DD45425C709F69982346E979E15C7ED5C616BC8E7CAE1DDBB6C400C31D218C8C69F3248FEB7D08EEA4FC81F143CBAF59371556B5CE5478F965F3C2734A12F0E106D267849C8E5158BB1D11FBBC11E96019B37FBB5810C7DDE0FEC47309CB54DEFA26620E89D79C807E8BD9B207C3C7E536D0CC53C22EEB39DA5D558BADF2BEC5354C2BF31AD82BA70C49F8D1076220EA43A8AEE37C34EED45C5E3FB7384D164C3701464A6219973F64E08EB799ADEFB7117D1843D3E0712C9604E7D380A59F2E8EA47F0764A009076C43B0017297F367B8836AA26B0907CC0B99FCD32856656A27088D329909A870A2607756394AB70DB9C49D4F2465453EF594B29986E76AB8E0E1998A81B05F70E73D698CBEF894A2AD2077059A3E0DA0422A1B4981C8D0D88391E135BFF722B515F054BD94FADEF3003E57D636B9FC15F33EFC3A955C79EB825B61C11B1E52B04E7288501CA19D80B81C8A3899242B22B6B0897899DF96DCE84357DFE09B87C5FF0C5D238B6F2A041945A58F929F7B9163CDF2C47797FAF093D3B91993DA38039547951693BDCCF20E23D686206D03E3D5FD94497C28F74C797B9BE490E71BBD4F7F6A172780FBAFC6899049AE9E3483BAFDB709D0D6CB887DC7F22A27B33A2E2C7461838DFDCCE9DC030B6547E21789805D6AA5DFAA868221844033B4268117AC84706BA0C8538BAE75FD2D36A7C652C58672C95D75FE6AE245EB33762DE1EFA50ECB7D9A29C02C1CE0B1A9292E767E8D3F1CB8ACAAF106ECD957CC2CFED1C11583F2D82632C26B4980ADD613AE4913E1ABC5117AED3F5C5161615F721083B80751AC836827BC90FF38016BF985B02A7342C0DBA5422B5B4E16390EEF8872A42DE3CAC9535F60402714085A4D4849EB67B49194A9FD20EA0D84332F5890AADA690F4031D26DF747FCEEEA58E14787EB6C7E4E00C52E4C4C126D6892E2DE3212F2E49AC83BC2B00F7EADE11B2658A527647D11EF9EB502554A17DADB2E7B16D0C8BA084AB5D1518C3C681EC3B30ED1307523318FEF160F9AB9B27D3224BA95C68D373CC4BDD3DAAD5F028ADD05A5163D66F539613DDF66F06B34305D12D4BD84A6E2F0E04BE9E32F6FD07A8963D416FBFABD600157B6D1FBFF5C871515E1F7A51B58C92A26EB7BF36C4ED4560B7D4F4234471131F9079235134ACB254F3517382DAE8C73CC530FA2E9597BCB29EC79FE063BC82DC0A3215CFEC6D79F8283094E6C3F4AE13F14BDEED81AED5BF00DB512DCB8701BA6DCD6FA3F8338302806D941A3E90643432211F2177FFEB36B2760EB9DDC35FA62DB50B935618D0AE3CF2006A3EBBB011A1A240777A10A4EAA278BDDC505FB6DBCA2DB5D02B7627F67D09DF532120ACE516E12F4548D86F4BD3B7B8A616368CA90C52A035C5DCB9E302AE02FB227A82117B65140E0393D8AA96D181A89A9CE62B24F0910602BFE38A33370AADB4ACE548D3D9955DEE6AC6BD4DFC9F7D8986ED7C30A61C10FE00A4F974731B7F2BDDC8F307DF18C85115B15EAFCF9610A0A983D15AF63C55983DB77180D01A4988BF49F0D13B90DA38452F01B9F6AE9315C0C85C35279E905285055DB954654D09B08F81D8734899E9BAAB02A4B3B026FC596676C76329BAB76B7D512C0B625E15E5DEBCC85738C603D46E1DA27FA7DB076410505245DC1BBA67A6F64C29AFF4F8D54F2674A90B8F8840589D4FF6D09ABCD47B1CB6B65AB53DA8AA0179A0C92049F6F805181C636D5A6F331591559B10DBACD05C1E4638B3C0EE273C5DE44470C79C394ACE8288A920EC6DD14E6208C8FD1E44589EC61FEC335B2EC9CF0269F8C231A5CF7E71050E03844C9BD0138406C8ABA55F94E77F39C9D6046D3B38C4B72525E66A985C6901B135D8A120EB4F0A07A3BBA4A52D4ACDA8524C447AE2BC3BFAE646E619B1E8A9E7504B975E450045BBB4F265E0819611144911A989D0309B0E42C70F85943C09930BFDCE2D59ACA7694A48DC1EE31CA51B024EDE4EC02C605E66A1E3053631DD9E6A7D205DE395BCE2793651E553F87CB27FB4493B590469BCF575EB8EF175D423073B836FB27FB8B20524B3A82404C101768B3AE74473E120F1AFF728153C3A3744A4D999C2CB62241C375CB51FBF85846ED4F2D8CC2DAFC190FEA7AD6BC1473574D9C2AC9BEEF76F007F38B6B37470F5510EEDBA0B197347712C24C48FFD258A2A453AE2188F28FF9E2F5C290FB2EEBA42DD008D9F9FC81A4F35E0A4E2AFD538AEFCF1C12B7519786451C24889D2AF6D686B0607BEF9D0CFE3CE2C22849C26ED643B98E2E4A840B052AD85653C1300EAF81640428A5BB3F61BF686EA43994EC5185A6F07E0DBC9B45882FAFBEF241483A6BAD2F0543C8CF0A7F4E06A091092628CB919A29E44044C3A8658334D85F4CAD1DF78422B094EFE7397BA3E82D8A5D638424CB093F9C8BBDB9F75C0ECF7B40DAF93FBC9DFF9A0773E5C36EB065543A243CCFA16CC6C72C0EF3221C21BF9B901C59B5C0EB4C9047F0896835917CDD7E519D950A0BDFD1258D4E6B63A550783558F265CDAD8A31D38F279B1671C19151D5337961254D141751D05893932C3F7CD5C880411966E3B55DB29782C1BE23F73422C76FB9AA92038CBF1A93CEBAA92C8FF0F6F389FAC94239A13FD31F03F6D2FC02E1EE33D70D90A1B8D07382D878FF07500221A2CBA116D5006B9AAE1F30E31AF19B048857A38471DCB9A1C0D7D8FF7DE2369930038F0D2E1D45DCF9E182F4456AD42C8A131E19A36D7682E149B906E6736E89E0AEEBED7E5D9AEA7B40DCE828DE7EB0B0C4B38813E1E6F78187373C6B8ACF9EC248A824240374F5263F21F47BD712E6774DA34CF8CD8481F6C7194CB9882B8C99856BE6E079C38617D0E8D8A498EED5312855765F398E43EC10F32DE10A7FD1C248FD29B5FE6D2D7FEEEF09A09DC54D6EB53C695E384548CA74CDB0571C27B78BFC21FAF338DDA2FB3604698323B25826FD9DCE1222B182D29E497149E2E317CFB850E6275AB2353074F7423786CFF9A5BF102EBE02DA69426F0397BEE389ABD3A3D0ED134436388C6FBF1C48F198B5FF9CFE7EA0D8DB2F214FFC930040A8D061A9062AFD34CA2492E47B2E9DE1FCB856371BEF2C91280936C50F1AB289031D0BCD2CC197E39DF376E0984A9AA7C7EBD481A38F766F7D9E61D59D5D1F10384A6E7C6898C8338E01514C4EB3FD4A63A44E2F8267ECB52AD03F81E8D1BE7ECF471B24751126253459718B93B56A1ACA9146FE99BBE57F0617DF7928B4932817D5EC84108C3D60381CE82B91EE2049D377434506F243D3ADE5A02E6765869CF1B56292A86A35D5BFB7CC22E76DE3B59807BE2DA98FC88DCBF86D0E1B4876C5BCA527EC661D4401B6C0C3D9A7BCD34B87135AFF5882E7E9113B406B1559886A809C65CDDFEBCB489365571DF90ED2085BB38AB9B2A293EB8A8B5023D4E298575B1D55D437838FAD5DE7AA13533FE453684AB1B6E19550C1F45B4A35E5054B8CF3A72590A70ADB9535191EC64F1BA7C75A7689A0C5220BD84A452A4C95B42D32033E248B0B5F56B0928C6EC48AADEE26CE4DB4A857328904A6E6D8DAE19F062D967F82018B8845BC3271A97C125392F0039022BE7F0981F445F658BBC2320FDE8D237E306A6744FDE28D2B71E0499A2B6AD62B8A507118209185DD571F0E73F823E27D588679C45455AE50C39FC1746515BF719F79E3A0B016895F2E800E4C4CB81D95B5F92BBE00EE0EB3A34D03932003DDCDBD110C45791A4C2CCB2E8910BBF467ED114E40C586A38AE5D9C6F9E70179372D5F9073A3811C7E4030A18B9145AA67500BBB481A25F007B673569563CAD574BF97A9908309014D1730E67BAB0A7F564828DC3F415C8BEBDB672E479FD1503BFCCE1BC6BC72AF44F67B34F81147AA2D555548D00B9FB5B3C3336FEF0C0A3CE1323928DDBA579B3CA282796E6A89F14CEAF50B6E15F14A585977EB99C118A74B62E5A081E91362C0849F9DFECDA21FF643E436E73850FF16B866E8D80368F152946070C567B5E643BF858777990BA6735C072EB2A3E05CE1A8032A48D11B439F786CF2EA57CFEF8E389138135131E74E9FC06A921B3685471F2597E898FBC5DE2B5192C1E8D715219076FB5D3D57F6A89FFC2854EDD57451C301920A8FD6507CA69F5450953DD2D92C793B4803A00356D86B2100680DCA8EC91F13F203D4115EA8D8AED22CB9CD24CDFA74B00D464227C1A2E936DFA00DD05E7DEEB3A4C87A8721BFE69FA0A426D5912ED919489B1217F006B8315E2E91F6B7C69628AD45D4929EB5C7AE430FE75CB4701B78F445BE7F36E58CA2DE1D2FB37F0660E288423D1731C913CFDDC080D0E07DC6E55A1E7E67516E83B9DE14ADC7AF423431D28AEAF0CF5A14E1F389FAD4E3D43167E624113D3D1C5F6DE14FE3750894A16DC3E1897F841794F7F4FCB07E51233D996E5267B3676BD37C1F1B4B44CAE158C9BB7A07EBF0F2974A7D431C230A926901DDB08F2CBDB471B2DD7F67F423BC337B9A9EF48CB4FE645F94207E9F3E44B535B93B46AB36480EC73FCA89F669364B3F4C44594C7129DC9F96AE83C8A4D88E625D1828A06C27B0047157C12F966A314B2789DBCFEEECE335BAD782EF99117B0B35A00400344F8894154EE2DCA5C5F04183B2E3A8AE812D647A2644C5592466009C0329B4690ED31B8675CC2220FE9A5C6E7CD527CCDAABA0349B5044F4605D9402A6191606C6AB54C72D6F16CF316F966B54C3CF250AAD837BDBE896D7FC7125837DFDC7D94A408C03BDB4CAD36B70400A1752DBB18F6D19A8D44DF487FE33045AD04A5EFD7FFC428A17DB3364163A7BFA2097AA957B205DD268AB333F5C158C8351E3E5C64FC172C8329677890BCE669D7A227677F9DFB3DD812C5FCE1630DCECBD0BB7F479AF24E7386DD07277FBD529272B37FFB147239E73A88D8D004D03D29EA4C8D6B2493C6D3ACE8AF9A45AEED9B468ECAF12DB318790EA91984670F1F98642BEB58A2F3B7845F7007B6C2C0E82CD30816F96FDC06BBDF1358057FCD042D94208D0E01590154E7C8CF325E7EB9EA4504A6FA77E09F8915958F7157A8103B786FD2BFBBFC09C54D9CDE01791D5BD9C956A9ED97939CA3730CBF88285BFBB4520201C5BF790794AA0B8BD4634AAC505ADBDE615DB0361A2CA1ECCF81E3DD286818B949831A54B1FE277639BBB60EC1D3694CFCADD310DBE5DBC136496AB927B5AA0E027D9E9C0A99FD19CD26CFD3BC00202675DC106C4110106856ACCFA90480EC56D93F7E7C378991C9DC70AA268311910E4DB58EC163B8079D606BCA68921F40C6FDB19738813588F29FDF1FDCF3B3944869FB165A6AEE5BD252383738FC916ACD3FBC96504A01D151B941F82EF6CA647A1EF90559E775DBE328BF166E9614D04D447628DBAF795E61F747E8758D0A0D413CD3E96B6DBD322BD20A6482A7ADEF2DA4FE03DAA38DE4790978650D1E908244A652230BE2C68E1BCAF0EC8C84F3942C23193DA9EB931AC6C6BEF0164DE46CF42176383A2AC030C8842E8DEC2F8123B2CEE941E160BE72AB74E5F3380C1EDDD1872C1FA74C8215DB0E7A00B3B01D12C42D4FE1873F09AF729527023070C76B2E2068F2C564AAA742B5B21D73F004E4DA586BC51750DA0284EC2D9C4FFBBF52BC8F2FFA9433B077D1A0190DA95A8BE6FCFCEE8C028E85414B358F5D447FC50EF83EA954FE398C40D62A494B0457921C25E18B218AD7583B34D648C964134BA064EBD7CF31A4FA7697EFA71DA8CD5B906373A20FCF066416571170FAEE4FB22E38CEB1A2F314A1B1BECEB1EC874EE2F811EE2BBCF7D4A378E1F18E1B4789A1E2D16C40741301BF75BDD9C65BFE9D8D242BCA8B29C4576A8C67808D652EA84CECDEDD6916728C978BF382F4E146897A21A74AA30EB9E7E703A3C47686BA47533B3DDB8BD402E4CA7D1B6985425BE1A4B82D0371C7C3D1023901A708BC4E655297AFB50891375AD57F9DB7B1B9C1873B66E6E7D028D6CAA6D6B1152DDEC4748A18246A009E9B707CC6A0937F7DC67F126D61BBB950A9629B9BFEB97A84DE877BB4D6618FA033C9CE505CDD5D11AAD14C15EB524C38EE30DC0EEFF493F69F847B0D4506DA3C91C88092FEDED7DAA6E714A31A0ED57F3F7964956CC93126AB1FF554288C03A82A5EAD9C4C29B157DA14C79AE172E3D8F581E38A7808412F3C7D59C345AA64EC2C05FB43B34576654A959371E1308EBDAD92BFB16549E224CAE9DF8E9864FF08AE2B8048CB70D365E86480B753FB23FCCE40DA5BD0077BBB62F3A6446445CF9DBAEF092E44485D87E7CCE3F37A84873C758524C643B8AA9723EEC723EAD60CC20F98E062609BA7E714E4B70BD574BBC0AA281F66B150D5FD73041D429F7E4D2F04A97BA8CB3898337018DDC93A674702BC161E25B7B43CA2BD65CA73F82742ABBB33C8E1D4944A75C8E52DAE3CC66D973A1B0B34B6E58F22BCC9D19A0756B66565664AAFA303F5775B5ABF2AB47B981DD25E689FB78315D8BE7E52597AC13305F28B59EBB7CEED95B82BD5EBCC994442A0A50F4D907410C775135F195AEF1A3B58EC9BD28FF343E05456F15EC4366786DFEFD6E390A992883180E89DD54C136B8615CE703223B726D05689A8C991712E5828175C3F3BBB0199C0A4B7BE01B5AED02157FE46AAE38AF7B080E6A5B0B05CF0159DCD64C124B40AAD083234C9E0846380CDEBDB45F8E53E99DCBFB417F56654C88BDB41C38115A27D782F26A09D6A38E51BD8BCDEEA045FCB083F204342B22FCC5063E69F4EB189837916B6A7A06C06246FF73ED45F3607AC1749916CF525B4100A5AC6313B9446EE63F603C6B5997DFA4FDD75EB97A2A8CD5EE8060DD38C8AD9B64F9749EFF2104774E19483CA1A5806D9C0EA9C71E77F1B95D99817ADAA5F837692AA3025DF3877D5869BA66E1C4E2E2C761291CE00ED6960DD9E237C7708C80459B3C8DF5710943B7F6BD3617832851EDD4CB830D30949C9FB731AC8B23E6BC442EC6319C0D89FCF9B9FBAF88C6BD7A30338BBA4DEEFE7CC3490DE7040499AF5A6FD595A2C35E867888348178269CA995F9AFAABE5A19A8C2C109D7EFF00B15A672DAC935D3A7C7D6A41B90C9BDCB5A434D0F3A87CC81D02AEEA0FBF2034E331B1DCE56AF0CBDD21A69E0FAD4D9712D9AD5DC3DEBE01C0B6A132A07E9F3EF367B171C9C79EC590D55F3E71385CB05BEAA79737AA0131DA2D65FBD02ABA733D398E52323B6CF9C03641CD9BA4040D5E2CE567E96844246702C74E2433FDA00AC1EE32AA09D4D19814D9B90A7A457D0F9636BEE24493366DB23BC0CA59FF7D2CF6B76F863D28E8EEB9C3C269C411A753C3368CC85BDF4E349FC374348F7047002B4E1CD3375EFD2932D0FC8F903527AC6E3F35494288B2B716B9A26A7BA9CD9AD880ED9C04587F5C0C6F53AE8C920207FD4B126FF05F0CDB481B925199C470A3131B16A32B764F20E6A6541049EB0507EA126E65C5482258BE8552F57FE68BA3C6298192B9670AF47B1CB134613FCD5AAE3E24D4B6F7782676E7580ED39D8EA75897C742512961FDCACAD42DECC73A8022A428B8A7D72E40E9428AC2C1C1477CCBE1901A74BB1978AC15A512A47D5D5A97162334AB095073664C87E62401FBCC96CF5AE02E3258E34619CCD27DFFBFD083F13F5997733932B2E5ABB32DE03AF413369E55AF50FDED4BEAA2C9E912F9EC0214679E32E3895096818A1094D12288E8B7C67F201E634CA30202492E12529D38B3DCD696B905AD8C6DB93ED2482A8E4E26AE505C16DA7513147D7B6D7BB8314A06C99A6D3872E8B89DC33F4C9779CABFC31F866A07EDA93B4176A0C03486CC67C2D0C8B02E4F12EB050C6E671BB14F8002878EC1C281738083C2D6589BDBA65879FFBA58A1D8568DD26D0ACB06AF65942E94A4C39AA1877493EAD3344E092D3FEF10DCC682E01F7E4C4C953B025246F84AD4B977C4D7648654931049C3B8EEEB168C40CFE1700EAC6346D72330DAE2D2AD0675AC899BDA2D3196F68BDD0DA6CB816E7A5FA968B24B89B63081721B9E0CA83523B385158BA0DC5A435202E91C27AC1CC8A2A07F071221A5476AD805FAEF8BDADB7B095B9059813CB39D8EF182BB0ED14F3444995D927C25E5066554329EF8E71E338A62CA2C35EC1B8C112C09AB3196B951C1FB50AD1292D077AE24AA63676793C87F13760A73594A2CDE174CE4CB953E5A51DFD4308472EC2E32E357337D50A9786446F625383F15408F567B1D8F3A306D9FBBDDE5BDE06C44B0EA13DF8885EAF23F0E9494E1726AF92BAC298A5722E79B7D5D6363D1ADFB1B67E0984DF61091248325D3111B075950D74E160524F4A8545797183C8CEA1EB9360E5BCC63E0902BFB609F5556D148A9CBA363F0A4568D725AB64F87CDAA14469C0801D11BCA07938389C4FFA198E75E66E287687499C6444D4729621BCC6139F79666A38D705406DC62B0A55CC573E0E01D1104FF8D00AB4A2EAE58F3B78544FDF5F3E7250B72F2D6B80CF13C4DAD6AED56138CCFC49DD2A7CBA60CBCDCC8459F58AFE486A0DA044B3E626448265F75922DA4FB0F7B5BB4CA898A04BB5B6F18DFF9989C425F4B40A1ABCC7CB52F1344AEA854CCE7E46EF2FCA026D2F862A4959447F9B8FC12A30D4F1643B9F826203E327B18B7DEFD1F06E13B06A93377410C221A32C7099EE5440BA145E61FF4A3479D5ECB5423C2C662425DE7AE7A961E826C4FA29F1ECE5BCD1F78BADA640D89F50AEB682078232FC30F1699B4A8A0635FD80FCF960E28ED64831B8849B18BAD8BD9E6E5B931FC95C34C8C8A1060466899381F3219906D379226710D9B28D00A5E5FD0C087F30988B40E996ED24DE24F2755015DDBD3BE3AF53041C603FF37AC94586866DF1169FF925AC503BB3C7412FB86484DBD6AD8D7D5F0F5F33271CF738BE755E0956158F9211B48E389E76C8BFED542265ACA5F6A28547C980E659B4AD30A7CF03CB98EADE42572573B7DBBD73EC1BD90523D8416BE9BF9CCFBA437AF603855EF0A348A4DF4F243E3597A911FFAFCD2E10328D3A9C893A8B0C3D12C7FC06DC20EC0D3DE4A652E7E19B14B6D5F8BB7A680F5D4D1D97D8E11A68F8ED3C6D35C4AE805BBE98D34F25C22CC2BC32B2E01B03B84B7EE96818F331BEBAA7F34B1372BABC6605EB5A39B5C0738C8ADE77D96130817F8AF416756EFC5E1224263B4E93E91C315A509A3D5CF61A04711478366AEA5BB625068D260723AB3949A58F5DB0C48F4B80773AC3BC5EC07F026A506A186CD8021C6422EC14E465F9134B30FF66B0EB5BF62D5634AFFD3AAD3A80FC3512799839C715684BD08CA5F5AE4C4FE85FB7BC35D2D6AA3361721FB9B7D3DF637B6C971189572DD5DBF38CF1FBE41225E6C1CC0E76A3BE17CCDD9D8A92E703E02C5A5C283B9F36308B17069334B4814E4502D09E1A8B4E5AFEFBD11D4A91526022CA89DFC88530D23E6CFCC525953D029878A36B5C8596F28C5CF4E7E82130574E5BD0745B69BAE2D721AEFA6A08E72F246358C86D6BE124C1D4491388F0CC5032D2FA6131212F9F7DC8A46A19487D956288B91F931BA7746340D4376AB2171874CB61DF20B1CF4D672F05063DCA384294BD95C37807ABC3115BB63A7C2EA58A4665719565AAF6A5EEBF2C91C8380ADAAAC2DF3C5A431943BA7453D5465F02879C99C58BBA2CCFA683280BA1EB98AE9F4F812EA0EC8D4DB0B26EF7F268B7EEA226D211EF535A38C77E491BB4DE34C31CCF10D13CB2685FC5D66A91B70ED1F1ADEA52801FAC5F5F9FD3991F4148348F9C179C72A626A906A90345819956B9A5F0698AF63D2DABEB6E3315F91E30FDC65D2B0931D5076BD1A575773BC303C958889D6669C34D936AB17D1D8F77DA48D822659FC2B765DF5A1823594887FD6657A6DA3CE7E5E83929D2AC288B67D5FAD7109AE6ABCB997B9E0F1F3E42DEFE05EBBE50D6EA5D9E1E8F2A7FE390B41485F798300A5EA322DE1A85DDFF0B8C11595E8E2B78978BFF0259B086080F0D690DD5DAA6A7EC69F5456EBA8222C95588F0DC7BCC098E1D5208D2578F889347C2546E2FE8D5D289D3F2BB2A4FDFCE8C973CCECFD21C280CE31EF20B3FC337A4BB0D5B1B86DC62C9B8970843D6391610AA31D8D99A73BC6C7662144EDEED00FA5B059FC22A2EE4498723138E8CEFB611F65A986F48F7D7C0E371785FA7161166FD607A681519F9A4E409B1BAEBB6EA2F8AB3CD4A24F1C1D436DCAA812F35ECACA5FFC8AC56A2026903DF0AC1E534C4BECD84EE0F41FA4C4371CE7648EB525C44ABE54A5765917BC1AC94D3A0241C21F7FB844963367EC47D83A691FF4CA5167F89AB1C70C351D2875B76D0B325B57B2B0DCE8BC6EEACFC95F1073F296DCE92728364B2CAB233696B153105D229748AED2969A0CA27B19CF8391C6641442902A73A1B77D46EB442228B5DC383E98788C02D822CB5C567E3A8FDD24C5290F0867C5F6BE1241C37D2D551466D54044F96756B089EEC350367DE96A829656F91761DC82B3A5E5A3B0A48B696888D44D4E408B74DED07EE803F7EA411967554680EA418A5A28739AE0C1D7A634793A107A2180B3A5F364164B9C7212A5F6D7A2E139B8E742690310D0F8D3D8447AC71B2C8222A8275B902C570D086DA6D009CCBA1B3826A12FBEF4BA189DF76A73A2CF264233A3058403DD96AE7F3241609435D4661190862BE47385B0C24CB62CC6F40A3498A17F02639AFDDAF3B6E701981488F2EAE8EE97072C9E7FA3A54A2835FB4030606DD65B39B8E651A33997800AA587E909A1951DB179EB48BE43D07E814C460E067E94D21A698F4777BCEA903455E4B4CB2D4503765D55EA711616C7B8639268EEF375865972C6DDEB857A8A02BBB75A946409E021236C45406548655DAE7954BD0FEF9AC406DD370379FCB15C26E848A4CA570B0D054207F511A13E8B7B480101A25B8D580243EBE9ACB240FACE369128629F6F55FE70820B687E93C5706D385A6378EA46142FFB4D6E5FBC77D8453783388305FAC980C1B0226BBD7FE5D7AB1494626B8A73DE03DB1BFFB84E5208457B7700FD4DB4BCDFCDCBC616B260284C654E4B1F6DAC81B28D01E8A5D70E27DE0808A7D47F3F605E89D6F70FD6F6F6E6A8E79714AB9C3FEE3CA914B1EB8711A3BEB717B44744B60D2F842693AAB22706D4F417DCD48D71B7D8630E71205C912107A169D74C3C8DABE93AAB5324D39B3E9641FA566F0C0482B7CC2F592AEF3D5CEB743B9DC0A39749F8C6449ABCE08840DBE42D6979F07CAF2CBDEE1E4F3CF08224DA548BE9A9737D05D7C0515B19269821C612B1ECA4C12CA8E455A862E67BF009EEEA851B0F9DCF1D49B4DF29F9515A6D43CDB4F8970003F843B1BB5CDE7F74B10D997FF2F8C022F00FD803CB44DA7AC678D8CA8C92AA7F8859F26F8274833340122A8736C1F29FB57629451CB996773B31A9E2301A4BCA100A3CBF5B751AD339774A4F074842503C3AC729B8A7D6B61E61087DB14C5B4EB7325D9457567DFED5CEBD7DA414769C113306A9022F9D0995C90C73C3BEA75B440CACB9D0F1A02B933F91BAF371B66EA56548084325E30A4D4B5E0F9BF3D82D9CD9633ED4B4B9A6AE76707080C319242D5FC6907CFA9E665EE66F9B5D163B1064B5558A9B09E76A2CC8B071713BC9E861611AA37ED9712E586F33E98B9BDEDCD13CBCE96EF69CEBC835C3C56C77CB3DF1CDC7323F58B9DCB79CD354B75DE786B8E2AB23D2F0AA0E1084E8FA708EF2CE38297E4922C63AAACF50ED5DA42B88322ED1042F3B6D45DB152B884D9E551D8796916FE700831822F8E797B2AA706056AFE71CAE9B049ABBA218777670ABA5106FE9BEAAD0B2D13C5609052E4F36E09FF7E3F527B84AAC08AF070450AA2147413008DCE243F62BDC8C5C54AD2751D4F1899C7C7601598AD04D6AFC97BEC19A0AABEBE05329A544CF9AE6ED58B8C65C3E255476EFB87CBF68D08FEF03156F795E9410CCD59B619973F89CEBDA0E4E9080179D913E9F668073A3F5D50BEAB9777FD646C7C958304BEC1BB5603D844D936FDFAF6C1FA385A10D097F312A7769D1A78E3816BA97ED642DCA1BE0C2F4227758F6CCFF841E51274535882B691591FFC320074F448F53206AFFF5CE933B2DE928F2C811D81A58B69BA814BE7D2C19D5ACBCCA6FD52DD0E187B3B216B7C629186C5FC33DE162302A259898A7FCEEED031D873FDFCC885C70D1978EE8D470B39E6AE14F82D53DD1824FC09F1D3CE17DC5FFAF1D833AE8E262D41F220C3DD0ED18F8E98582B92292BE84AB7885584CBA99907B1381DEF8D0D2F1BEA766714712BC4E29584B561AD65B7F4ED9CA5C64B186751E6E9AB6DC914389B6815163C5961D458A470BBBA10912FB1E6DE482565583D287A3FEC7083857D222E04A76D303A38B4D163F47557A6E6E3CF338D1FA433C66CF84EB472E536BDB2C6553C9F2E4E25517F9DDB2A1D311690C7BFEE6D86E96562BA1B77776ED3301FAC2C068FE6881621A56660F961F60B71EBF3AE36A51B4D44E97E740EB192F796C7849B0A8556419516650B003C35705885A29535AD89408A9A2B1773B24BFC317DD8732A0A065636861C9CC7F507F280384C8C7D76EB935B773DE99D631E0AB48F9144EDAFEE654A1ABC4C88B19FC6ED53EEED7ECF098B3A8885D2407EB497AF31015BE75EEDAC209F080FC3A8CDEFD43B776FA78AE8716F5FFE66A64641E01BF88D18B45AB590C69D17C88B46361062BA71587F19B11D009425DED08ADEB48B488255E202103FD32913467F87DA51CE83EC855FFF726D172709F10E1D286CAEF85034E4EFD749C3C2C2DB91FF0767A7C0A71BE15F6ABF1B0E0762DD0529360E650CCC105A65C3CCA668D5A98399DCB29373305DF939742B0352CBAF4F74033E0A9B702B67623F8CB9A72D27696601D7FD5E66DCB8BEE7158FFE74F9FF2F49A03EDF4B8377F214E3FD89541420F651AB259C50654FBED2062FC4098EEC617C86D3B3781B42F3107E2E323348B22CF2464F9E802F2FEF6916D448AF5EF2A156BF6EAB3170BB257E74AD0228BB70960E44C96661B84959C0F273D55F0F5EE5D6C172C20C20C7DEBC2F7964033F2BE060FF75F2F6A81E83A6E7899F06C2E33B59478D78E077AF0EA6614136738619B29A5F9DFAD52A79C86087F10D1FBED8B47139D6DC6276B229CAD11A69B8815735C1A08671230D063A52176AA977A0C83B77A526B84A2A4E9E9EE56EF9DFC11B3746A9C948D009301E113523BAF99CB7BD353CD7531893E06EBF661C54073427C1F0CA49D08188655D0293AF2CCF88632D6225123BD0BA4BEC51D565D9A928FCAA9C7D1F3B3DBEBCD6325143303B9A5D6D98C36554143E4E82CB29423314389E6461DC682A4BB5E184727CBE9876541997A62FB859A8AA3156B7F8B1B4C1A7FBCBB3F9046B10775A163F47FBE659ED61EA26DE2FB08210148CA19D9B89DA126D8826A1DF364820F75782A68DC7B5FA1F5CDB8548CD08AE40B58DC5066B84F423F63C469E3F55547C6B99ABFD022CFE9D6F5227082A30CD7DF876F6C9258CB0A37C97E4A8AAC28E80E980AB6C549A280A3B487BE75157D246E7C9FE0B1F2530E0A4226274AD5CE43317D07FCE6CDE6736DDEE8DF8D46BACDFD42045439E14F16A480FF31494C6A2B29C8A25B5FAAE3D2F61FF71F2C9C4893A5C81FEBA0FF3D656EE2827DB3426D889B8A88AAD21ED0A21AD752C203526C65BAE5977FAED19B0FCCA3F0E92ACBD45F0F1B3BD7FBA0E74782CC80D8BD90E1770D779E7766328685C235BA122367A1F5E725B9E3D27E7AFD94C8CF42EB6A12FAEA433C585C2B8E83B955C8D170A31EC2D02486EF62F223C33126E6AD6DBD5B682589261A0183F568913F0C384799421E386985CD9B96DA4B5C59573A81E51FC60C410434AAD5ECFC3C5E1FF879C021E9DBE24E782CBDAA27FE899D9B362DDE38323E65EC1181FB3EC0D1B743E53AE5655278E21BF0381CD23F1A82E075C914C4CF68128213BA48A2AD9A178DF2604580F4D7FCA960D2D76126F6E6E1C373059DE3C30B2C140C0AAE4343C1E65D2A4C4862F204C92E3DB1DC55EA9467EF798B3CA4C46A50AB55B5CBEA567C08C46C84A2E14D2FE208718053277EC54583ECAE2197D4035A2F55C2DD1E4323F35ABFD15F01CC7D3E9DE407453EE8EC1C229AA42D09A9E2A8B4A124FFF0D98F61C674110D99ADDFEF831D2E6945BA262FB63D2BD035DC47AC6C6BF751ABDD6DC3E055ED493FF3E63B880D03E1464317058464BC500E2AF7CEE386766A632398B736423522CA590098240FE1EB1AC9A3E90396FEE6FA344BCB2D66B49A2B6AA3250670317C8358369E26816EE19F15F9BAEB72E12B102CC21CC992C80C30805C5253421F35C18A339ED6E4F7367DDAD01AF398616EA2DD53F41C71295CEB89B4DF1BD9366F0FB7657FDF29E46E1004D86B96F81352F1636E10F8B172907B05F7F0B7037CACF255E95417986FED2934D7FB9E79E987AD8A417DC2E066EC2CEC38226B498A7363FD7ADB506DCEEB73541804039016C1D4623A17448A9D01AF0CB1C5DD0E270263416B23EE66DE787029CCC386EA0DBC47BF3190DB4E1F6FE199206AB569E55450335228F61C92ECE09173A475DEBF3A3948878BEF03416725CB947CAD835466D62D45A681CDD50A575D62059AF94A0313F32D103C6EEE64BAB4A428B087014C45065D836E9C59DE1D10CB68E69E4B9D97AF0A88A114BD3C63F333B9D26871AF878183FA18EC9FC8A166C9DEDBC67EDD9551FAECA48BF5B5BD297877EBBB5A7D496C49B7D48FB906CCC0048344FF8B4196F51CFD9A251AE429C63178678408B74EE85CF503AE95D761C2038A5863CFA73B35953C4392CAD8DF6F69324E747A64559F4E688E64A3F8BD95C785A52CBA8C2FDC1D07A8F7E7240F49EE683732C93850DE792D0DA545ED2F3E6B7ECEE8D7E15FFB31A07B94B466C9808DC499FB2FAB5B49F402E0EB4CAFE721A7BF4D7E0E4416CA76DCFC896437755160B65DA0EB383C2AD6C26BAC2EFB0017EB5BCC2A9E7DC9A4EA2D92EBB0F9BA011E04D3A2D511C26B93F1145ABFA96005FCA2E50F5D1162AFF23C7CD53BF36E966B233F8C88A1799156BD8251BDD977ED23C720646C53F2E92E9B618CDC48520C36AA374BCA7EDE7DDCBBE51959129C824C43404A5F1A859BC11649FEC9EFBFE1EBD2D7B41E5BE6DF2E9B5E812FFA662712EEEF62FFF3306E7A677CDF3E46291BC43C85B3E7762D1CDFCC96885C5008FE63EE2BAB2AC115ACED2FC1281E67B78FF58D509361C1EBB612D1C81648B16548D74AA341AFA452DBE4F7B6713E065A8ADE699464A4351F979732A8BCE9C47236E0B762DBED8D9C2B8DF6B21E0E745F2A8032B094DDBE13B76BD377C3205EEE8CAFA36408AF979BA72764552DF523245BE50FBF9B2661FFB5BD77001FD6CABC7FC45A01B2EF73622F3AA66881F2B3066BF33479CAE52090C8E7783E4112A9973C52E8DD775EB806E11F9B582ED3D563D1046912C80681B3C70C78508779047FC7FB4A9415CB164B9F40B8E429460B9E2ECA4176226C4DD24AF13535C3333714D71FB9D1EBCBD77A5D96BDAD819E81813C90976A5F265082598191B84FD83D8BBA69620A273E585A927ACD7C51617C37E68E6C5FC5A436BD978AA4A0EA35395F9B915A88C1B346020D369CFF527A8A3B4C47B7A8E46907B5B55DBFBDC750C778E4CFF0E1F04795E36027E424B872618C517C12DA5FA5327F173100E545F8E150950C7FFA737C951E3F8F60CDD897F6A014495563E80E896442905B81400204C8B66641F083F5C5FFC2BA04F8A32D6890DADFC8102CC65CE1D6CF0255B7426FE64801AF50F264A9C6064AE75652B6CDE6F42E6CA7AFA47444A0DCB0DB2543943FFBEED9BC97824EA8D694D3C3D82E9467AFC5BBCEF70D8596334C57D70E0B000E339BFBC94C5EBD28D36B000122AAAE0C380B43A7CCBB044D8773DC004186F785C69332E7DEA3D56D450B5E33609922A84700C0FFD304419878BACAD19ADFD9D5CA2F4C7A49B001FF6DCD7372BEAA5BE7F5A01997D31FFE1812135756C947C9E2D040DC5C0D60CDEB5B6F8BED6563FB7A06C499A9F41379B6DFBCAE0015046BD3461F9514740C5F5B24F828B0A8D84437239FE92F19DB12C04BAA6EB4048B1544E4E7E022CA0D81E904373A2A0BD7129A8366DE3F8D693C55920585133FFD8DF9C9B7AC8B285A51C0CC65071953F08E0D54BB0DD8F906679B69B1C0E823EDAFA929255892257C4A5D9023EB27C0D4B09DD245C24493ACF5D431804108DB9CB0F5B3BC711A869E6D1662D1535C70C56448F5EEA12405ADD2CB46A9D30F5A166A161073600D0328CEEFC4F0BA6137DA8E576C8968ECE54FC31D129E2A336F0338F63D74BB6B440F0689B4FFB136256A4D4B08B4E0EF4DF93EFEFFD2CCEF8338BD7A5F41677D30BC3CDC6A048F84709E4F5B0CA8174683DF0D841D4215EBAB6424CF9D8F7CCC79CCCBFA915C1269831E0EA1521F95CE9B28D7F30C2BF1591D46B3FBF7227F5C8C8C2BD7312EF4294BD748758130223CA5DA64DFE9812168505E510B631D1FBF6CE596DE0A8D23FDDB8C49DECEBE87E3DC88872E30A9BDDDDDB38AE6EC3B7FCA67A4497CCFE24E4D2DDF867F739F05F16A9BAF46F5DC3D146C4D580DA10A0BFDC03E7CAAC7D537BFC9209FDD6EFB04977B52563422CF948340AE8661740A73590A9E0A3DD51F771223BA12B40BC9C5E1A707BFE254E37747230FAA7EC2265BBB8CD3DA9B725593B1890C66DFB2233F65CB13E6AACEB3B82DF6E99F66C86944A61CD2F1EC573F606F0BC329021A706164C5914D6AC51810E99BF6B1B8C9C72EB2A5E0EE7FA8F3E95472A08632B82B23FB883DDE99EDBDDE382F5DC9E9586245AC3D62EF0E6DC7DF8D8535E1C94F2127FEB8B2BF009D976622FE1C6620E43C4EE983AF8147E9D451BD7DF621C037EC2F08637F9C20DFBE9AF3D62BF260132EE11F41F7CCFD189A7A7DBF01E5D0038CCF5A3365F570EE97D77D03A3FF772A8D05ECE2F5B7E3019E8B060BC656A34BB7C968C132EA140EAAE66A7E35585A0FE2BCAA8C4FB8BC3D537D64F0080288984BF6FA8D33579889EED32334B9B929C833F13C8090B52E2AF973918AF7D83D2380763DBE2C29D27F0EC35352A900F4378F6E6B8AAA17C59CCDC274374C112AF9F446E877AC8FA575D7982211C013098E033069346B826018AA6403EF40D83A4F9C1F99A24E0C26FF09285A89A85B28007C9A504CECD1AE7FEBF3AE608A1091F9E7E26A58CCA60B40C73834B65F130C1D3BA6825EC726038873578562221489ECE773D8566E43D5B91CEC8CC7B5E6E7BE0B78D87FB17F921AD3291331A9B98EF733DA33AAD45872BFA68D4B5994177BD7CCEDDEB1B68612C64118894CC164185D62E3D88B6EE52AC559E1BCDD61F9037F9DE829DE5FB9782FEFDBFEF57DBB09AE8F139FAB39745A4871D8402AD417A97373B108F94C91EE936C3C900A5A7F182CEAE5E5641E68222979C1DE065FC4C283B049D748B8F2D8CCECF883B15E00ACC7C3BADF80BA71CBF26B762C60F6DAEC262C002EEAA412D25171123C9887C2F486503377A30700083A4FF1F837A2521479B4A811EC4D543FFF379E4E141DCA41567989CB6433C106D41FBBC65F3AD4859089A0B1776008C7834F9A233C6443C04875DF6BDD3A5062662074C0B334EB3807D34CD5CC9A5A3B02FD95C1F20271B8CDA5F8FCCC44123CE6A3C0923271BBCD4023010F29B026EF766197EA8B67DAB691AD471E944094C08C528FA086E689382BCB21CF5249DBEC2F3C1C89CF6ED0458561CCA09A530C4AB00212810139B3CC4F408EB895B0807CAFEA84F4CC7168BE3092B59A7A54F72D6766B8138CEBC8D52DCE37D7079E119BEC59FC6F8F7E13C68996FEBC4FFF6AB43A2B32A267ACD71A03B0CB74C9A8C25BEF950CF585B20595D4E5F11DD6F6778BF002DF331D0D46893155A53790155111FC11850A4A0B62BCB96030E3BFB6F818FB448E1A3238F3EF738FBBC69A66796B477D647AA9CDED73AF2475DA5A2E504DD42378706CEA3CED1EE8EC1A2E4E1F6D2086A5E14A0AE5E7939CD1D44823BF95407594C94ECDECFFBBDAE702B18E73575384C09B84FE8095994C79ED4E740D80B673037B28AD2FB6CC7B7154558AF663051B3B912983A5089A7B06CF847E56B25632608C73A35D6E9EFE3EBBF91CB8BCDF8FD14694F7EE6EF1E94F657120451CF0E54BADEDE8FEA1A02F84FCCB11020E77F0A0E4DF632FFFFCD99503C1CD716D116780BD1DCDD11A8BE156D4DF04B41F6497318041B1BC2FC47FFCEFBC587A5543DB6E2A89CE0D80D17935A32E39FB60936E6E3943559FE56F05157815C10571A2BEC80F67A809CFA2047B4FB83D4519D46F820D000E5FBFB4A844BFEAE7D4121E39ADF09583C57857B76C778BDC6A8CD1DE1EABE66EF29A8CA6209D2E685E2B88023700AC0D4AEDABBA44C7D9FB406F1687C709E3E86123E0C3A2551AC9A0E5394CD324B39C992162E2CF62D70DCCCEC3E32D2523EA6FFE2CD4491F2EDB67F1C265C47C59B69C20F2CD80687BA71B75D73DCF4FC3634E3B6AD3F1633D7CF235027408CBE91BC6130F2596C0DE00CDD94E3539DD25A98982E461FB41792083D90665737F296D2B9B2E606AA9BF53A67DE1E41D28F179E048144FD730B5FDDABEC2EE86865E5547454E00161D719862BCE125D8AFC94397DDE43C2D52F0DB45A9B05220C243E25A1FCB72C3545DBDE497F2771312492B56814D4B81990A501C1E3B529323473D618CE036F956E0CA1D82F5B37C6B9068BBDDBC483E33CF3E58D03619A71F9DAC88AF343E507208CD3C8C4B42B7DECD4CC3FE128C12ECC9C162874E6A4C4A28167FEB8D418614F5BB209ADC12DD24B4F446452F4B2ED350E980612ACEB2F93DF32948F18860255E8354007CA481F0D874314B10D77D1D719CCF98C6D9F428B6CB7899AFFF1C6AD4A0CC9C5C1F1EEF6451BD0F1F9EAE76B1771D253A1F9465CE3E7C6F1E52FBAB1F1A45611A599944437D8159E33962C3BEC49A5629CBC020DDB78251C288989B26B5221832B470266582FB7E24D2445BA73900B18744EE3EE6F3EDB9B79C7CC72CE32D0AAB1C6F6C2F22381078F8B5AC1E4D9F60907F67FB1A714BFB0A67EBF9F8B6F6939C8C8C5B76A99BC691CB1055003AF7751AFE73DE51EA3E98A3546A4995342ADE92551A21D94A03CE9D69FC6BC1DEB8BC7B8E25A578AD333DD2CC273AD9A2A3E9F233F28D3FDC4CEE2A211F6865EBBEB479372AD4DCE46D5E2D2CDBEEB8FEC4F1AC6F0E4ADF7EB2FAE82E7778410AC77F014008A6A9D88450295260EBB84453402F2F2873F698E9DAF651F32C6FDE527853275F86467696B581D7DC895042C39E65B6D390C94139F519E2ACD61AB34F60FCEFCDA03D63F6DA9F48F816F9F4A5D350263DB882A7BE7C4F6FB22388AD654FCA9B44BF3B2D1B29CBE5B31508B5BA0A1D1337982E78654BF4C7593949C043440B39F8BC09BCDD5203AC8536296C32C9875C95F6F149837165879C07FAC97AB765836C84AC4913F4CB425FD700B4B07B827B3F8F8E730F4C487A4C23207B8BCFE2C8B6B3E4E6634C41C7A520DA3F39852B334AE52E64E1664792197867146B7AA438D1862A3D38AEA70F80643E5513FB9B95885E9FC908DFAB1EFD3B11B1D6EDB96B9B9D6598691DB5FB2DE5D30529DEF926BF07A2FAEA90BF08F9455FD33294EBA427C0F1186DE9B719A05F26BEBCEA38D17E26096705CE1E0DC9079B052377B078F5963A72DB0F4A6D550104256721EC57265749B5210AF7066C77C7673281C58D90D6FC3E5A54D4F8834D1E9CA6B74BC2C212365D90318D88601E5B1188AB3EA6BE70865745BDD0AC768B55CC50358A7C389ACCB133490204A8D693D37370AD1A10F05F15108C735EB5C78B98408186252EFD479109A29D3F460F0EFDC87D42A00C5481490B592C37F8E2A53CE742A705D313AD568FE067EEAE171725E7E24F1D8C02BDFF535CF622F76A21D56E18E6538C6F0FDB9CDD2262D836F2E2AA801618BCB93CB04240F778153A2C4161C2F380E88D4978AEE24E505EB987819AB22D3D687C13776473E8DF3617D282A78CC7F8D4BB6AEF7CACB35C89A707CFD12E82C3931E12CD6DF0A7C10BE7A608B8CF5420A171B5ACA5944EAE0EFF05AA262E37AB72A2341A87DF9F13E702E666A30584A12895D3C769FE619A47B9DBC060AEF4A13744504019336C5BFD7E7996735143CC3EE37E73BA49B6FAB9AEA45117B2E9849310846734CA1E20E543BE4181C84237FB8228B9595126B7BB144AC9A43319F820EC2A074D1D472279FE172EF55759D588782053BD1B2FCAEF9D6132D35B8B718E36FCA2AB8E77492409AF1BCA1FDD363DC3348AD492F6A0D024FB4E9C24BC3DC3F968B12D6E6962253E05251F7179955B829BC8EB4961F20401BC6CC74E3E61FDF1693D3CC1FF77E50A02F71BC10113FE68B4C1510619869AD5186ADDABA2848507123832D26AB0A0C34AA01339DD2330FA3FFF1AB680DD2BA9C1F2D0E76533E7390125C3CCE3FDE76B8467943BBBD9C68E31F88CA327CABF7FF81F23EA7D55DDB60C8B005AFA3501A6273A0E46F078B985B12667414BA347E644BB49503CCEFCE1274F36C5BE67334894E37249DDD62471FABC46D9F5C7ECB95C32F37ED0B67BCB42660C985D758E6962867AF7BC6575E9CE52C2A7F300F61FD571D4B63B2BC23B9263A79DE023659CA5296C5C5DAA240EE90471630161AC1CAF895E0F648CFDE22B3BA93D0F4424A1E02A781C81629DD4BBD4A92D61AD0B347B9639F63038712BFBAFEF87CEB513A7B3BF03126A8D0DEAF3652E0B0D6556E6EEA8E2E9997B5A132299D1AA0F26A0CEEA835EE23D5C63A681DAA1FCFF00DD819FA98D9AA50A1CA027A2710B829940C00E9C3917BA79C4E68F432EA5AF5C2AA0E86DBF170EA32438EB559E0C93C52C269EE127AFF942F5720BECA5826995F721FD31605B5BCDF18221F35B934F229AC598298301BF5E8D70730AFA60C5CF217D7223131B210F5843A798BF3E37A6F82C6A530D18C8D4414EB09096447A5F2EF68E2C54EDCEBD8FD72BD7452A521C332CADF3A7080CDE50C55695A937257E873AA6630895EE4714306ED34F7BD424D7710F83907DCA7CD85D844FD5E8825A0497806115343C852DE6BBCE31D377D24D26CBCA2DC4E43550C23E3ED010539D67F2CB6013230985543262AB5CC9E267070684E333FB1FF6906F5AC4AEE518FB8CB9040AB648747BD31B44D5A7D892C14D25E4E1623E530F4655FC11CD58A195E3BF295EF5103D2DAC6F33861245606E37C824B10276CE234F8F3C332B4F6FBB3A94C45CD8742D98F67757B871B17BA972B2F59874AE8D71B88B67CBA735D7938BEFE90B5A318F421F4785DA05494B3791FF67E96C3E941FD77FD0C678EDB8B77445BE2093CD856A887A357D49C8F4720B1560BC4324EF993DA4ED8586D4EC1CC9A9695B9067CA63374BD873C57607F09029B1638913FEAFCE690D9D684EC2764150653FA2EB0EE47255CE1F800FA664C755158F68325D7C1B71CBDF97FAEEEB6891B8BB916F14FF1780A1414922046F26CFB97DE33E1B7225AB8208A40741DA8F7E8EF4FB5CEA738AA5CBA8C56D62E0515D0A1F8661CB288AF006FF196F190CA26B91BD54EEE3F29F1A64A2C96F93F40FBED1C77CA86941321201E2F360BAB259F0BB2DE140F90EAFE58AC448AFE91C9691B4EE5E42674B361C6EE0ED798B6470DC6EA375E2EC679F4A17C84BE28ADB471F8B6F8CB6F06E54A6D1E9F4AF659ACF9A6E6CBC9999EA3E717D3D13B87B6F2E7D8D5E7FF3C0168EE437FF6F196939A377C4F2FD865A3864C62A137C7E62A1F3741D79B3619C054B9324F7B0FD2E1465F752D8DD4131FC6E2BF9BEF4F73CECA6C19C57D0AD7AA7D3701DCDA86C7DAFBAE2C2533A2DB080466EB10C91C6D9CF35C2FE9B867AFEE5555476D7195F184AA2FA80D940C34948CE2CAF8B017CF99B5A5371FE87BD97383090269D89EA89F1E28823572D901022DF9E2C800E8EF3F440260AB1F61D3842241543A4C634BA3AE2760A5E1260EEBA79CE2216B1F31166CC19AD1443C5D0519BCD173BB36AE0F9CB64B4B5AD6AF9950A736E69744CB863EB718C0A14F31C3F8A7D5B06ABD21AE38DBA43A731016D8E082D6FD473B7F6C18223406D39A7B7FD0479DD43466B31AF13A1E028D3B404BB441891410A5334BB9ED80C92D3922AFA59C6A88CE36ACD9B6FB548A2B0949B59B185EDCD93485930827C7C8C9C871ADF35FB62D5DF76EA922D82ED91435CD5208A43590EBC8C667EEA63BD5C29BFEA0CB532D17AFF3AAD56668077D56FA45B67F236D65705E09509DA27375190971513CA4E570C9C6F2F8CE52F53079EDAC95C653656ECDBF05A28771436FC0844C952EFECFF24F89EAC03D2ACAD7C10F14996BF89944C53AA1D73EECFCDE14049CAB0D0506CCC201B520ECAE2EB459D3724768145BBE5770514D7503A95A60444A918645754961E7D223E779F21A98FA99E4392473426937414927ACF166B5197ED2DBF3912A9035A54DA245EA6F94128455DE2DF6527E7796812EFCED819691C003A4B8E4ED340C9359B9F1CF8CC36E14F85433176573B0CC106A872B9F0BA60846BC8977BF906346C5E4D7D0CA2F7FBFF3D82FFAC22B4A6D0230719D12D4A4C54C321F961DBE55F67667CE58A88F1729AA126E167883C73DC95F65C2206C0CE9FFAC7746B3A0159959C64CF7929930915DC542E329D4D6080A8110AF906BF15E40510919E2CBFC2462A1361EBA4A6A3DD18C918D85A1928E2AB34D46F24FF5EC895A4BBC034353184FBBEC8BE0352392C653D494AEC049777B49ED6DDAF54B664D5A5CD6E63A2D263DDE2BC5476307EC27F69C6D0A91B2CDEE9BC9F731FE88B48A841A2FDD56EFC8CBE57439F8BFE86D7F44EFDD13D5EC16C9272C99ECE396A506D3DDB6A889BF7A507500CD6F477187378C346E2CD421DDC79DE335070AE24C4BB3ECF70E6CB100B6A5995663EB51AE7062062165DD438140A43890B2A791E1ED6723C0B8FB071126205B7B1BB60637574D2FDDEF6E4CA3AFB93A955937B035C0AD82EEF56DBEB7697154192B1E9F0B932AFCDC171E345A801938053E9E9EEBD5409CC26DF920F269A84E8824548494E69791C99D8A31A9EB04519D11FCBA603E07593375CB1836FE189E98207DF993AC842368D6DC4EFA667862EB42FE4E3274BAC4D604FC0E45315DDF31FE8CF86C2BF230BF4DAB0348514C22BA2B7973619AB16BA8568F996A1C09DDE801056312DD0E78E474E452A65E99EFED3D5AA74019F7DC2DDB01E91987D675C215D83E23CA8D6630A9EBD3570A487A6B1467247AFC509B6B35167F38739C4E19F2F7E7F40B827CD094BCEDE0888161EB6EED97FC9120F3F1F016B239EABCD37515D7B27A31239B8855CC2BD4B28830A896E555F1772C7B8033365D2486120217A4A2346D5A233ED112969FEE1A2821E07B0A2D3E79E3BA04D3F8B4543D09E0767829A623C44F302548F2B295154BF72DE771FC54576A4A9BBF9D335A607E494E455C403E17753DC12FC8B4ECE8AA326798E2BC44DE3B548D84D4CCA3AE3D28673A5FE7D46DA0A382BE4DCA62EC188DB83878B9EE09A93002A97869947D77F9D93405232188642B18CB740623FA6058646675DFB1C78BA1B215718DDEC13A6114744B8958F4EC24CBE00C8B7C4325FFF323A3C9D7C6E3293A8A33A9990A2B49C2E5D24516FC519DF78CD15E459115B995E69F23A67012530C3DA891110DC9DD89F42689D043391908E255FE2E878DFA4187F63E6DAB2D79914BB0CF5BCE664182632DF69D507EE596B011DABF270384DB36396678F02F9E4BF756C7AFD2636A17A20E24CD024436FCE3D9E674D40B232CA43635592937A1A4C5D7B94FCC4E377130F73DFB78EDE0D0178E9C5FDCD90EE973ED708C4FFEB39051B04711FC4442A3B17C43ACB857DDEE21475592C03DF894849F3563328D8ADF8C06E7C68E11BFD772EBA7CBD09B32E6D23473B02E64F6059E3384CA01C1A5129E84842F778B3422BE06BBD9EF30B5BBB3B686DA4B43DBD7701C4778AABACF9EA91EF2C0B8703F4D6B0F7083C7854CC7DB6312CFC5E06AE8E807E2E2B2D3E4EE5EBAA3C70BF60CCCC7A54076E6637BAB193F8CC7CB5C5A6911D48AF5A60ED837D6934F1A713E4D52FB5BA81DCC6722636028B969DD1480445F0D6DF52BA504B5E4D05A664A417BB37A5C41EAE5544E0FDE59B8B73CE48FFC3686B9969861774676D34AB35FF9D957682B7BF8DCBF1005A5F1CB24A0582394C66949527B3B9A271EE1EA9005B7F13EBF80A81A1AB74194630F7F2AFC55428047F4C4221B3DF25E7AAA55B2394CDFC604D4F4E99D2D5075960138655F20E780EA24E6350CB096ACA1A94AC705A6C0A3B83271EA744F1E96182791238D7BE990A5131F5B9B6EEF49E20CB5905B610B665EE8C768CC59E0CB43AB68EEF60FA0DB19E3CC1258161D0061D98EF8F686D22EE6DB550DE78F417470D0C03472DCD3C27AE50AE17EDAD9E1C99300267DF8B53BA63578F9E3453F2EAEC3906CF8FEACC6C11246A483658D16509FC27725680EF553B761DBAFD29C8A055506B276570C3DEA6B88412F4932ABEDEA263554B3A5DFC419A01B618769208A5304D7E0DDBC466971B40B2E624A9095643F7E448456B37EE73B5EDAA77C49EBA71426F26164E6C51FC0CC91CA645960DA3A79D3AEB9BD22C27486D9B865B5505D2F50A8E2FEFA24A8DCDE4911B66F95391FD4A7489465FC2083EE4246C994C04491C839FC1D1181FDA31158BE48A697D960F4224E46765F43DC8A35C9687E18EA4D82DBC0A6CD5B7C29FE4E1FE1EC8EE9B82495A2E4A3D8ADBA9F80C3FC05D5D83B91618F814729387185500A5F2A27F7E67680AFFA25967D23B5DF5383B0DFDE25253A2999A057BD478725B47D9165F7B2F1B17E6C63ED60516DBA01F61FA4C387637CE517268C717941583EB80940413ACC25AA6BF07CB3795A40D42BD4FC21EDCE0870B8AE9AB06C72D2CDBE5876B80ACC03C991A486E3CD22412071CC962FD6AB38061E60DCE68F489D5620CC94F29DDA2F4C2F1ACCED162122FDD435B80D1C3568A1B918CEF10589DEEE83DFE5F9AC897B7214572494D417C93088A22730656A00652622F52001443ED47E8681D1951B1D8F695EAB2F3B9BF9C4B91EC2688D48EB7DF4759FBF120F406580AD34136487692CB19F95CBC2134CB47EB61872FC340F09BC23F9FF678D1961DA56896DA1FB030C9569ADC39A06D6262F5EEAC129BA6318D51D67960F334A67C120800CF9BD2FC4C20029F195002BF8C428761AC49270F18416058EEED6C5070EEC750A2C32776515364037DE85D54F68DD2A608253051F1E895F5818C69C37C0A829BAB7BC57AA9EEA243F5D3D29832789CA5EE1C9EE83808734D3550A3631912EF456AE92A69A710ADA571815D54D32B495867A254AD53CA1CDB28AA1680E414CB4F5C0794E0D49A1E3EEF40846CEB778DB589A2E7460D397541DEEBF4909298D2C52817C2BDB8C4D88DFAB01D5549C13AA51E7B20494F823FF77B2A88C037A592ED83FC7FCDD5BB4495F88D917BE4D2F02E419429301BD727B10BE299816D82FB3D2EBAF9C4AC032384AAC3E758E4B6C0419A5D3D97919F5C3176202B1F31A39F89FA14781DA6AF83ABDED2AE54E0FEE9D0B748A6A51520CA1E70B8899ED194F222A789BE7A3C072C0248BDABF9DA965D8D339E88CF43891666096CA7BE87BBD0EC6B0D3D619D8D79F8389EBA203A65F0C0201A6713E713FFFB24ADF64351A30653984BA4E6B33952F41BD314F7A00668767EE87C63F927A2A53D8C7533AF8F5A0D16C85445E782D37F2EE880E6EBC36A6FB715FD4A19DA71F968A4DE7CB0F5B53C0A210BFE3EC47DE10BD02B99A7BD49728D90FDD1B7C78DCA6E25DD61DE7BC40F46A2C3A13527B6707F46068C53E27DE1E44BF9BCF55AE2E8C2BB9E2EFB98F885668C170801B0877FD9BF41313CEBF05E5D22D3B4C025573FEE105B7B9F4F41031B1574903D5E3674CDD0962E21EEFA74F81C433AC75A6FF17435A96CF10A234C0B84966AECBC98F43C2FBC83993714F979B2284F968B7E9754FC0DB9ECB65880D0272D200591659F12F2BBD0D84BF0C3988836E6B4CE69747B413D940A8B90B6B26612308F02080AE22FE6DA4454E78C710F97C54270038DA261A60F3929A7131C5886F01C765852CC36E5E414235BF73E2A6B456A9C0AFD8D7DB488E7796A0F7AC5CB22523524AF794E74822AFA991CDD6AE96A62BF9510037F19FDF1802174A3C43E61A55FD9E21DC0F4F51D70CA305B36AE00169FD88A3DCF1AE184D0BF4C3B62D301617038D8523409ACCF0C46FCC377F82CF749F57F8870DA3AD9F94FA3F49BD1AFDC1ACF6CEEF8E36B14796E10C8F6B866137AB80813AA69CB098E1929B80FB6E3AAFA5F79A584E95F4AE588076F7927AA0976573B67E8871A9C9CEB7F54A7B9B2B3800123E8060946383BC4B37570454F7A38466F08028784E30AE532769FBAC00F3E26A02A41F8826FCB66666F1A16F33021F49D4A82972F5D275912D20E714CBA16795720696E733E85660E4E6B833928A3BE5A0AEBC443B595EA9D570D5FF9B8822251C0892EFFD1D4626E9CCA617AF9080BD3FB951E1BB927207B48351EA8131A91E3A250EB63AE77EC86CDEB80B5ED7A4946639457320C6FAEDB9B6739D9E894082FA3674C9063017D3C99391C4D4C51002D106D7C932D29FF83FE1EBA1878DB94DA1D20C7B0F51BEC37B759B8D48E684686BD720BAFEBA231D2506A52CF74049BD39D3CF165AB8B9C39F0B21DF4D460439A9FD86AC414DF9CD759B7B910298777287D8486741310936D4505ED15019015F68C0C16799C34B755B63F18BC35EBE597A1047A05945FAEC171F8ECD0B423F9607A0A2D3C153BC7508C66295B0619F952AF68DC6C66A23F5B9440E21E4ECF8E028A24D14769B53B39EE1DA4E9C3752BB286657334DC49FAB07A6B704E59856DA1CCC9C1B6045FFB4B0ED7E8B739E3AADFD0A6AA8E94342F45212C46B3F31E4494EF28CA8B2C0B6E244F8DB78ACC398DB3D0C2401DB9473B65EE2B77851B6B4DBFDC675A2003DA5DE5A652FE0FE3A40751E59189F0F15554DAD78F6AA0F52797D9C0A2D783AE104B4273F50451EA749C98D2B27783549E73BF58D1B4A1B21EC4DB0096E6D8E8C1475C27CCEF7FA850A294E95131CA8C89358FB23E680BDA1026AC299BB043D7394C0A38D87ABE78ED2980234AABBDFBBD946F6632EDBD508EB964CC1596C4DCCFC65A1AD302A41CCEA79038E008708033B51072FFFC804C30E5B9CDE98505070A27690CA2A27F2B9E57A272A2032766C8BFC55A3BB9E638B5DDB946474DA3FB707BD8AFE0020C968BDA519020120963524FB84A3A76E4EA2F26F27ACD31AA0041B079FD0935FB847980EC1EEDBC4A78A1F9263E353DE5A4C574BA613B359370274834747496B5FD36DC5D68B9193FC9E8F24272FA79317B2C82A9DD9BA413E3BE6358180D9A5E8A9E1547D54B5608D5607D8D9198E92833EA18DE201CB0F814B63319E5FD8358AD6FFA071274902B65BDCEB65A7331373FA0FDF21752D97699579F87F0A320B19BD8F2A6D901B3B4EB544988A2A54009E98CBF6BF0075BEF9399DF4674A02B5138467BEBF07F26CC9F56742C9A20E344E7BF5876A84D2F663CCA813A56CD7D6D58EB350B8E17449C7653AB8D20792B3CA4823E7DF12ED4527EA685A457644742042464AA684E51E352B0F94C65E66FF82104E68E21BF415CEDB6F0CACE50BD04609934A4CC7E39BEAD6078EA01B37293BCE46D1B06F9E903A5C6E5599475990B7813DF186D86377A8CF56F9E47C7765B39A87186162F8CF7A29C43465413FAFEF0EA454DA8F58F3AEBC7580F890242BF8793B964EC9913CC94343A466537769CE26E18D7DB7646C86D802911E1FE96F3B53DF506B963566AAA34890BF22E209294DF9E56AAD772B34DABBC63D6F9541A22438DE41FEA503E4B0155788474CB3F2910571488DFA07100EDF1915E315FCBEE4081E5093EF168CDEF1CA4A93DFF23F81BBC9E107B334CEE97AC279A4BEDEA3644F25BFD29B12894CA631CF0A8BF7D3FD2940022A443E76E8520310A2E2C968C993AA49866D9977D8625E90AB3D4F4B7CA4664446EB11E94C2AB92512593BD9475B22C5AB458815456D47490FD837126BAD9802FAD0B7977EF1D9F7532D4AD9F4DE3803A049CCEFC01B0C48FC62D8C30B35B83C18CD5DEB55077E4FA9EBCB123FF53A8A8443B4DD09A8B02E9C970DB995706CA345A0927A5BE60166934635F9EF441994AD54B3C96932B84995B003D90824141CE49B4B0795B495D3E2A96A333DB972AB16773AF8BFB2125E3D532FDE228B0325690E40724961E7B29D33F822D6DFAA2B30159481AFA1E60A2F3A8E26BC7732BA4EE9C9322E1FBD334437FCD9D3A67AB22512E336D24E89D0E7DB20B0F9C60E04297E3F6E00DC2E4638690BE91D66BD6297E3E3EE335408521FA10EC6B4CBABAF71A7D32FD2E9DD80A968B91DB9CC103D958CFB243D343217767FCA4122C25E5EC9492274D26A31C7C0057340BCD9E0F5E1B95890487D50A422FFDF4C14D2F55EB3C727E87D10359A70312ED6755CED34082D26ADE7FF36F45BCE63DC9EA9524B142F60C6E03605A0A548FA798F2FF98629A7030464CAAA153BDED2A0A64FC7888AAE3928329E5731739B08817E1CEEE060279F4ADC12B452A8F21DCFDED785C535A92EB4DA17F861B72BFE2F6A319DCB85D34E834F2B6A40D9516925CA070741D8C1AAF7C79AA58F0CE8FF17D16E11DC2887FF8F0CD2675B494BAD122B88E445730D16C4686F38D985EE33CA09C0A451175BBA245B0766041AA8A055BA0D20E872319F6B23153FDFA01B72BC0070D8F75E91655FC29D5971030F63AE10F602AF899A746B88EA5DD9B251A87E0F2D2EB4C9F4805DDC8E2D86AD90423971F3EC8365B6C2BD87CB78BFBEC80A0CF500B5473A88F16B9A4E53851EEB23C7DAB55D65A1BFF6D7E2EEEE993F7A451BCD2EE0910F57C37439710CC650FE6855DE6595BE21157A0C729FB3DC1F528D38B5FCE09A72CB4B7DE3E57D9DB6E3A1DBAE714566121903B8CD96CCF0FA583EACC597B333729C5CFF2B4C87F1F9664FE107820259B46416061537715E769867A48AA6E758CDE7DE964A2225031FCD1F7AD04E1F2D6FB4F8286337E4F1AA86EC516E125483DB308EB4888CF275C4C088DDB1BC950A9F6FB8D8FB05447BCFE32D062A1F397489AC1824E82E329949D9E52B6A6A399AA79CB466E946A3E89A00AC44E4B7657E065E4622B416BD67C3F15A637D54A7655735E58E12EE57F305B2B5E9B7AAE6F71B6A10047D903D880438A34026F369A4C5659FD706472330053BED45C219A813C22C663E96E6A39E8455A121E72E094E0C7DC33EE4FFE3B9CC152C6A3119C6A393F723526C3A2D804B5CEF8BD6ABA3D4269D3C64B3EE4A72C97BCF5329431E6128CD07ECCC4FBAB6A8C6D0EBA60AD59A5C49C8D5C227356F3584A7B8A6300D42EE4814CA61A923AF0AEF05566A4F0D39A029ACFC3CD9F1FB1E24867A223FFDE3B416FF44F68756AC92C09C7BA15F54FCF0DCCCC6FCC2E8A51ECD4879BD43B672E754AB2456523996605F68EE6306ADE84A0A58AA7FABDE703219ADBA7FE11E75D9725131C1E7DB0234482EAE8DD6FD1BFD64DE8D136A4C2A7FAB002832A290A7504A7536C5CA70B1D307EB1091347A31DF66E10C67E9C520D4E555ED457B727ED4B3D3E75BC31021DDD5720B88A46F6EC3C6796B10EAE86ED8C4A5A44570E8EAF0D29F1BD0D1F4C91E507FE8534DF1621973A2F6A783AAA78C0B5EB4DD574FC0E5C9E45F913EA54BD09E707FDB358EEE91C44EDE55F8A52824217099647DFAD23A9BC38D55E7C844EC2216F09270A80131983EDC887D16683D3A03150ADD08F3608A690DB739C8FD123A4B76A75A2B98B35A4A8300B1EBB379C97483605AC67AF9827DEB8C4E830EDF05B575F9F10E74C98CE60603E76448FD62E1B4F128BDFBA62F9AEE43BC88ACEE4F39CA7AEC0038F012169F156364BF191DEED5D3DE6897178FACDF74E2834C8D5B1E1B2080E1CECD29CEBE89FC56BE5049BEA36E668EF534ACCF6161E89D46DBE71D52DC1F3A75EE41597C6625910BC96AF9917EAD12E9F69D9528E28D917F3E0C8A6B132C2BCDBD1AB927A524B6F2C8FE33D647CA0C31C43B2356A649CC1C83A3FF48BCD49721DCFD9D02FEADE33C689C02427634766E090F91CC2A6A449F3EA959D5980F58EFB609698D76F35C9DD74129969E3BEE3323468FC93BE66B1D66D7EC4410A5D6A1CFE1D66B71756E87F0DD0190289E5AC20BA91F51DC75275859BC8FCA50C0C67134614C8DA5AA418198BEDA7AB43AB1294E3EE7D6276FD1298FA812D344634646CD72CB834F87931F674487EBDB8D955637B002BD9F9CE351B1FB98CDB3936C582B37EAADFF8D510CC22D10B56253A3D1969EB046770F82E4F42ADE26FFF1927ECBE0E731BF09A1A17C92527B79AA245273711DFD7BAF38EFB6211F38BB17266382CD8E04929E18F238238EE234AD0EF55BB4DC83EEA28A8EBFA58B06D95172616E0DDFA4EF441B2CAC9180DB9C6DDCA9BC21BC5E0F59A1F961D9D749E6CA0E0CFA81B444A1175AD7D2F37F01C5B4D7467D83AA6DC126E814C3EC739CABFE88DD8ED580AF77B280293145505D6067C6C0B45AED1B8630212A76B0498BA4805D44F0ECC116703F26E530BAE55E746EE177343C383061E7D397D183CBEC6AA3C08CE52BDB03C2DDB0B732C9D384AF98A8B39396E3A0FB71D9AFB7DEADD233BBD3FADD5D25C87F5FBF8DB65B72CE5F7DB3F1358F1765F655D38D3F6C4EFFAA9D82EE8740EC0A4B7B4D69A9042523FB5A214C2772637CE1F8C8313E37B18D9C0BE9AAAF67988F4C6B75E22102EA6EA5799D052AA7885E410D2C315D5ED60293DEE245EA684187AAC6819A6961062A840CED774726F842DCD75A7F24292D25335A764131DF683E6FA0B13751BED77E3823C2C5ACEBAF4D2583CD649DC1E407EF9AD0BB3D757435F330233EB099FDC58D85CCCAC0C955C37BF5EBCE982EEC3BD1C793F0D35C1B7B2ABF9FB671D6DF3AD28DF28B95838E477181ED224F6B4D1274009D5393BFD7C19ADF1A9012D451AB94A0C18F5EE146E088DA948B8D613D2467AD60EDE9DA74101D084130D9CCBBC0060C5EE6B5B1CFAE8D721B69CA9A87FFAEEDB0F7629A95B794598EF8B63C33DB901DD99BB74CF38625F3935237CA7EF34971B663F651544AB7F421B9339CC398C3D42A6FDDFBF61C1A41EF07E0760DF4BA94B973D80E309FC13F31443CE9FD238494375253F8BA19FA8C4B89A7691C408A3AB29E463E50064E46D2D0AEEEEA8E4EF4221689DAE2541C396BEE441537022A0E64F624D8689F406D507F8DC4A0072273AD92A2AA245EEBAD799A1B1F549B403631D8648554FBFEFC97AE700198A8B654A5D6C32C426BBA48CD9BE0B3FA84A7EE82A96D9478BFC41240695CA44B1C23FC4E9D42DD39E27FBCF395B52FA98176095895F9E269DC0438BC5D6F51EC1CE85EBE2023D2EC8664D2497762E05F7E065DA562DF272561328ED052355EBBE1BAA5772E7BFE48392DE59DC6BC10BCE92CED866228003F8133FB5BB8144D4F14CFE90017DDF51B84E87C0BB2133CBA00A1A51775CBE82307B35B3FCC34DB577BA275017C929E45A9919BB025535927CAE8BB9590601E1237CD86BA2D9D3BCB23B7BBBFFB7458187DF386B3E6CAA338132AD19D547DBDBA0563BD9E3C8D9267084857584F0DD09260748F12064E89A4A18D79902385D9AEAFB671D7765108ACBAEC6FDA2CE54FF7A7D618A0C8C13D0B60F8B0CF014B79F2EEFD02422E1A7C51C13CD3DB8A42F014178676E2CEAB18D7276D46BA014401DCC029ED1CFBF19EB4FB15542CE5CE39431FA5BFD8E0E306BE27AAC22F534145137CDBA81164059484BDBE422EC6B193F1C1BE2C4FE6C1BEBC1C5F08790CC5A1323D2FA41215B1AA1734171BFB714B89AB9F061BE15796017C5AA5AD7C67F1214AE75D8AE0C5DACEE9CF6B02042A5611233813B9829C803E12BEC91D521052A26575A69D5ED3A9838C502976C83D499AD3D1BA30BE42D93385B5CEDF2C265200B096BB19C5F6CD52261D6F1A74C47B6787CF1AB184D951E8FE8F4A40FC1E46A68C5648DE8300FC46F51943F15840F60145047114B366E5147AF99266E0DEE0F3B554467CA1C14713DC66DFE7452F3342BAF6C10B23200D51101744093D262DB7A8D4A65DF14C3913F864CD050887BD7F8FB6EC91D81EB501FCC21BC9EB8B2622D89DFD075678B343A97ADEA166358B5B8991298AB8F2D6D6C3B1DAECDE0168FEFB7347ADE11AA7C5070683902B61D18E8E7BA5709E94915800CB05CB99EC7A849F682F7497073BDA70D66CED15C7E336F840628695F235935107007F940994A78EB1683F13AF91CCB926EDCA52B86EC3CFF154F46A77D7014AB1EC945264FF6342A469C022ACD075C18AA7264B3CDCFE140DFF7ECD7CCBED98C6FA2E4397F87EAAF8AFC51D24F9B3E71F61C32389162FF7D45697BBAEE6E05CA5DA68D0075E2947E4948C2088EE77C124476B5173B6E835DCF4BCBCB48B021B850522208D49F68E6A090E19535A08A1B560EF8EBF456B529DDEEBC98A757D9FFD30F9B622329A910B900ADE190C84CC144F12829D4AD252965AC21853672D5B5D9343AF48704AE1A429938F996444EB2C6F08E3991101D7269CAFFFE50B93BAF75A399A2C9476C15CCF3D72105C9E47CACB3DB267B9E2A9F9AAE6DABCEA3CACBB454BD7B36A08BB18830DE75E2139E82F7258B5D15660E70FD1C8201C3E0F939E6FDD8627C8A32E33F216C9E0F473D8860DCD934A1534CC91FF9C5B42EC3E811DDAB22253E71377BDD9A6135CAA911939B06886C7CE16D76B1BFDDECCBE1A895E45A92113BB92382915C6240642E07A639E693E69C58A96BBE6FC03E757BEFBD14D6DE8BF5B9148C06D322334407782FFBC763E665777945BBD5F31A5623BD64ACA282E21D1C96A54954294C197491A37DCBF9DE1BA1567645EE9ADDA4549A884D753DCED5EED6FF96821679D02910C58684E045BC14FD175245AD59EE9B9677064D09ACFA505BC87822821C9F3E5EA84C2B7002B790046613BA805BD479049923CB0FD705485823DC00A71FB580D4D49674AA560C75DD6E987C7BFAD0A6A6D6923C21A4C514BF189BC43672BF3BE20768EC780B91AD6AE633D99C194A3AA6E8AB73891DCD8E65A9D3639B34458C5DC1FAA4BFA89C6D0C124A12D5F1A505F57282F4FC67B7109BAA7BDFD463B859D1B3CAC8E79179056E8DA926984C0B50E9E78C6BEE811DCCD1647FDF20A3933699BCC2431F36178ACD3F5AC172DB1AA43DE783BE926402639EB48B9965C427931E758343425873EDB001676E26F50E8C869C48EC48FB56515B4891E052F3D0523D0F0F5E66D21D02D60415EA5332CC4EFCF9D82C0E5C8210F58B1651CA7CC0F4483FD9EBF54AE117D51AE67C0615977F1532CBD49E8BB917767B23439EB666E0F75272B4C0B9690A71FA82522602DC1E26572B9FEDE3E15B81869F9742BB37D4F1825555FB2955FC211B135727CDF24DF634064C38872E2B0A4CFC344B23A5A75AC283D9E35713C6922EB94E9ED0D0B6061D9A1B253AC2D10C49096AD26EB9E2AF518F1805A0C554E74A882C7C9F084B84EEF45BC91F33BA9EABD31DBDD9A7EEDAAD02A513E8023A5A765C9C6AE2D91690023DF76D07DA65D8D7F198FC00A73CB300B4EE50C6999CB367FC16FBC5183C4BDC2BA353FA047AF9D71F464BD69CF711BC8315484186A4D7EC0F3A5C49491F5D7ACB5BF801FD1B47C5779587B4C38E7D3848438658E00A6183705DF0CFC58C40BB4863223EE1F19203DE5A8904AF054CDF611ADB52147869E44C40AD7D3D6EC1238A150D3CC2BBBF951ED572816A5E8E6B203277A35868A6C1A99363688684E238D50E5EE8ED77E2737894EBFFE4019908B2BA03E4D57B9D6328F52882329D7BF1971A1359E2E5109B8C58EA90CEF5FF5A6A94857DC26AE22156CFE2EC0CE81135B9D91994A2A7D7DE5FC0376321BDD18F457C9FE2A2786F1758722656EF999B425B290C7FA85EE238CB7D3BF77BC23575339C32B4DE92BD0725CF24C39AAF30F4CC94EF600926A1D6AC2B2BA82C4ED6569D0B79641216AAC70905813CDFC0E870E2628996B359F7D85EB68397A5B4D992E613449CB20AA4E0B973A664B32E31ACD4EAE513F51FC4014724F8517DDEF13B59FA91DA039E6FE21DB4F9BBA6C57947C760AE189A730BE92E95620F09F8981FDBB688CB82447276376BF28F8E865F9022C57C32DD8570D07807B3DD36046DB0944CF7D509A28765FD1E430EE0DAD70DEB5096A8CB058FC03397A6473DEB1C066EAE760CBB7773B034EC227E861576F7E01C56AB4C1BBA6EDFB00C2763629E949E8CE02310D97BBA79D29A9B32E02B4BD6D8B39A21ABB20DD94DDF92E7395252A2D103EB7CE7073A1A90909F238E52D98B08446C39C26333874E74655AA4CD0C91A8D1399937656922705584C340EB2EF2CB3DAC7F6E98BA2CED15F47F52407A2FF323455E2A244B8EFD1F2024BB8D3B12867D3EBC7BC4DD1730FD5061A767BCE727893885313C72063A0B3A9E46DDAD21052C29C91B08EF29618E66AE58631410D9A90F39E62B53400BF7312281DFD058DFC0FE787E457121C14A08AB51A9E3B71F3E2F643167EC90C1A3CAB3671C709C86781587BD7ADE2765A980F3FC3F57D79F523037FADB4A81340960FE16D5C24776C8702065DDD69A03CBE8C28310B83FB0EED6A60E36442EB0965884CBB37844BEAB25937941DF60EEA004A54C1BB09EE528996FEEA7F9EF135253C31A19A612FCB6BFA3629A456592F150A7C650A48D1AFB60C18E38961211DA633AABBD3E54E7A11C3CCEDF67D1764DA88ABE55081D81B60C7C4386AD2BC551187D0FCA69FCFC54D6FD8C59BF6050CFC1329093D6B66CA856F791BF23696EB993DCB14478471862884823F37FA8A6206475BD5A90F2750DAA91F6BFCA57573B1C7CD9866B9FD368BFEE5737257143C5A768B87A7D0225AD9BC342D84815268371EED6550737ABB41AF1D96B903AB28F65E2FC4A221B69188ADE8EA6745D4EC3781031B1D8D5C7895D60191A884929AA059B595A3C96676275771A2484DD52201A6F0D26DAAA50D332A2E6B6D3BB93F1F6CDD7D5E3267FFDC9FA3EC97A0B9AA17ED8F99C094A310B3BFD763A294361DEFBC9C1E450CAB60860BAA8A7C76E2488E25C981F7459AB91689D7D38D6D24A3346A927DC81E4DF2E72D680A520EF61DF81AD6B7E528A7C5674E0014EBFBA5101DF88FA2E408CC1E1CF01592258A295C54B37787E91021F9675FDF580148DE6F9A689FD7C79645BAEA911AF80453B35D8ECE1CDCB041C3F1D70903AD72D9176418DD9142F4F1AC52528357938D0195083E0557E73A6D3EF071F97218F6FE29110A7584477CC162848C6162C9328F0D4188A48ACC397D3CC7185C720F9DCFA64F79D4CA6E2108C9E577372BEBE798005D536FBCB5905A3D6B4B9DC2459CA3BAB22836C361B70A3BEB91C6487CDBD7116B531E66143D3416B370C3173090463C93E9E55E8B598FF3C29B01E4B37A8EC14E9E0B7B3FE1364B71A534060BC71DE2313A3D9FCF3797EF69C5551D9E0C2076346CC6BC94E01BD5C9D2DA329FCA2B35155CF5B0E8BFFBA44D15FA46DB0E13B94A9E998AF95E6E83832BE7C59C3B7251328D617B8CC508B8A6DEC6AE84B1AAB4919D5FC8257A7BC3B8CEDD6E10DE6832D89B621034C1368854875AF75982A978B4D45CF80E60F67B755E6440740BEE50D2ABAFA6B422AE1A7336218B7C2D5C9E103B272B2277A1521A801F0B1BDE789B15EAD3C1EDDF7F8779DFB15A611E2582C4107CF6ED3F158E0EC7AECD8F02F97E6B74B0793C09424394FB1CBC0039443E00A8994EDEDCFB36F304333B37028A4399217F7E7E25603E8E0DD91A1A5574999D0F9D5DD59920BA747883F902E35779CC2C77CA23491B7CDAFDD0C184088B3C489E967682F88B17A2F083DDA8885FC2094A7304ECCBB2853E81A4E4E9D1241504A5E0F81FBDF4E3CE8F64B03A37F8BA810DB7C5DB44EA20F8AB251214DCD87307DEC014687055EA287C9064E5697127985632577FFBB17B805172F8C8B0C7D855ADDCA94B9208787F1D8C7410628FF3C561693987E95F758A183B01E64049A8B51C296309E5CADE2F0089ADF7F06833D25CCF226E8523668A57B2656491DF815EB00C7A4404C3F7B961707C7AC23C6E3875A9F59A0A3C4E8C0133200F911FB6CF49F7966891142FD9F6841DD8B54ED395D13EEC32226FF7EAF1BC3CF84243B932A44A52331194E47AD2B0DEA8BEBEFE410009D080BE236E1F7CAD94C6513C50D2F65F1AE4C53EC99FC3CB8D4FAAF8C0BBF97C69475B8757DEC1A772FF78B2623DE3B7DA1874F9E8E338C2E8D9F9E49B1150AC78EE888CB0C960EC156FF4AB3E4F4FE07E0B836B61490D702DF5D36A0911960D80DDB1CF6A31DD51BD6250D455BC11C3B20A8B8053E27AA163F9D47AD94767FC61A79869A75465FAFAEE4A84342B0D4AFAF9F246BAC95CE399CD82164D5CBA314B4E4650F069926649EB9B646221F34E59DA62B4E65BCB7BBB5CD931B6255880621FA2BEB279ACCFE46D8923E965972ED2C4AED722B23C869F0BED4FCD44F17AF69E8BD134338D7769846883056DA3F9FA9F0609358E5C133BE8D25E37A9832AFF76CF9162DE6E3731B0C56A3914AA592C8F7D9214706C72872124868D5894A4AF98871E21999851F39C7F016949C0304C80E03301F70D4DD18C1C5030A10A87278EBE7B3B003822B87D09AEEDCC2DB8F35E28B4D7B77C68DF9E0F412EBC005C42EB6D5FCBE5F99E34276E43469D3FCD216A99ED3E666AE4F1B38874FE15DBE9601D85E5AF63EAB8464DC18147C052C7BB3FF73DA90D74B7105FEEFA4C6BA58ACDFF124117BD9E12447D47889414B03E3F571A82DA0113189AFF78D17A2C41893DA774862369AACE978CE7D5B68AF79612B607654366AC8164421061E571D52722CA2203426454C07F2C9FBD74E0B47018DA1A1834B443A284D142D7A82F8A245A776C0AA1DF6D448533D0365D25D3CE2A97AC4421B958B3D12A79666B761061026A6CE847A1B6A9B9F84950A7A07F36AA9E722811D8BB911A09BC05BCF6C3592D3A8D44CE73A2489248753731B2C323EE55F24420493E830CAC453FEB434F442096A5E19D8FA314ECC197D3A11F69144963C64024F17A3C67AA7A390094732DAAEA9A98BE8BD2E2A6E5A09A232726E4002A91EFD58E2421FE2B9A30C902DE7E562DEE695766F3632B1FE007F646FB3042E13962602933E215AB68FBCF122FF0AF744D522942B7012760FDA1BC8C82AC72A721BCD874231150C60AB734508D802E43F3CC878274812C5076688BE7A963D567292E777A2FD0D39930BC02ACDDEBF337B37DA3E28CE4B5778F1DB7639D52F42C4DCBEAB73EAE1B70F30536FDF72BF8FEA9A667D750724DD1002D33B49DBC3C6A89DB165F14169190306497B9D6B0B08B1A4CFF4560E0F4F44B99CD11E903084E958136E05F4A8554D6CB0322CCDE4C730CC2EAA7CC4A361667EAE330FE3864C312B76A16B9373668CBE787E414F641F25E55C08EA372149F06534EF1541E01AF87A7A5D2E40EA3B4BF025C850D586290F698CB84A59FF050564D2758770363EB6C56DD794EFF4EC37434DBDE3EE302708ADF164C5C5B0FA606452730D6FE2897EBFB9A94517D99DF36431E5C3D78E34929FC4EBE5CAE08F388F8FF402E6CD49AD4AFEE70FB5A4A7AB45F5F29D2496AB90AB83C56641E47F1DCE83A84FA3018E065D27B667D5077979597643B78F0174C5A9DCF5DADE7226BD8D5E2B2ED92B09BC0ECAC3CFA7B07A2BE6F9B43E935292DC29AF89D0A63C68F8C47C9C5932497D27232E8BD734A3F2365D9855B63ABF158878CEC925D906889E3560C1873C61488CD8165ABDE2A11C2990A9E22E9E92B81B1967E3D64881CFB4BE6655F10294841A2FEFF3386EE75CF7646E848033DA9CBD155CAB9971B7346F5DBDB96F9189E507F8DE7EA85F9FCA1F286CE4BFE7B81C1F375A7B84F848EEA8D29211DCE18B70A7EDAB305BC50ADD79519A93D4F0CDCF7B09E643D5BBAE600220F509EFEECFAD08867EF860E4F44D8A9D20AE0F133404FDE7A5B1D982473775CB4CDBD129E9D91B29258F738072CF8407BBE131404963D9EFE629168F6113F942A8A1AAAFB105E6E0D80DFBCFC94D3EC8132845F1CA7B2CF0F4B12C35F09EB06A3B9E5099258B1105A7FD2BB987CA73C785CE6FF88EF42BA4320F93F93018C83C371012DFFB05DA442F91AD9E6891CE705E382DDF6D91A6559D1B2DB878DEF32D587ACA89C2CE6435035EF56EAB0D824AB5C82E3D30037A1E794CB4D3CA69FD6AAA987B6DD911DE6FF7DFA52DEF81266C69F6A4E09F6D06F7409FAA343D55C5CE8A34A84D9991C41200E9022C43EEB87FA537EAA068C929C08D35FA6F5D0FF3622349C3C91D6000337BCF5F5DC72FAEDB55DE5987E1CC67A3DAAC2E9C06313982952545D1F6B2F76AEC92E35733E31843E4C2C02167BC452DAF3CED9B336CBC5073BBC90F677436D50E15979BC89FB4CDD07E834202A6C4C97C8752C326D12C42F3736C7B487A268D81E005C1020ECA5C7B39C8993DCAEF3D636F98C9993694B9102AB9564107C0BF9823D4E5D90C6EA53E86870AD9E5642514843851D85F68E2EA6BD2E555A85C17AE3C0417B66F06EC9DE67B44B9ABD5C2CFA444223CFDB7E76FCE8AF5492754FA08897139BD8DD756C2528245386DEFCB65CE0AB8843231508C092F943557385429A6EDA9E08F81931BF918981F80E7CE672E612185099D94D805F25076B4C64BC2F26F880581247BCE8F36A15A60A7FAC63BD0F7AFEABA2FDD68A17F7111A07AF2A6FCA1B2C972D11B03DD5B0078F728221FBAFE925D54D7454E91CEEDCECF96EFED27572EF883FB618743F63AC022FC24BE90C718104A7DA097B2ABCBE84E99F17A759947616A8B2695CB9B643C01271329BC50808CDD40648AAFEBB8583435DCDADEB8D5FDA242A0C6CFCDA71FA7DD576678F3B46B5A107F120A9DD8B2927F5A913B0CBDDAE0AE0B03FCC0EFD8E24F299E5AD3CFB4E61E73F70AF0E0567520727E412D37FC2CF3DD9CD66062C417C9F5522D9F4FCF8B320B4770D1A12FD262046F4750D9BD1C91FEA17304C2D3CD562085052123C61A2F7252C5ABF38A43F314FA2CBDF6CC0B9C639D8CF7D8829877E1B7498CE7ED6C4870F9FA6FD407441EB6AE9FC1C924CA561274272C6E4EE5103CE3522AF5EE5D9357B1080949A1DFB953F147D866157BD96576943B8241A8C070C7D854070963D3872E93712503D37B4C0EBA1F19B6618F01055B5FA2C40A2799F7EC6F13D77D43EAED07DB1AEEDF9290DCBAFB10A7F7DBF231D85C2A466B0C98B8631078F5D14D8B62B312AA00FE91FA9D7834F5DEDD3D65BF1B5A260FD7F24F2FBAAA84BE2D6FAD6E55C9EE38EAD82684D766476CC0E53C33499716A69908C52238E926A0FEC4202B797FA82D8C0BDD093E8EBC4A47B5A59D7E9419B054DB0C5E57CC38BF8C229FF1FE38ED5DD9BB7FA3183E0E248ED04D6DD9387E47A03C26BDA56A7BAD17FC5165A5C5A0532C4CB79EF7171792D7D5B7EEE56720AC28919BEC8CCAE54DEB93F25D4213070E06B6C8A53AEA2F579A65048DE943FDD7512512B89E717CBFAB77FFD949BAF4FC2B0216E7D983646A8734B94E8335C40BDF202EC5AD04AF8413D6BE22557A4FA37F03C49818A30845D00EBBB7A1BA62EBCD089F44DDE622EA6D8D39AFAFD8C39E1A3E718F8AEB92845622FC7124B2C69C72CB6B80B6B92B8BE65F85F57D33E402C51C87A3CDA0FC82581EDCE67B913ADEEDD5CD0B7165581F64D8E9577B5D5F3B9FAF5567901D35FF4B557F20197A5F36178078C6CA92ED1E47A84356B47CB6420EB622F29FE78C5C2A536C10276F1E88E15A29923875E94975231C6AC57703FCF77D11D199A00D1AEDC7B06F8E5CEBF02E330DD6C7D39BA5E56FCA56F88CFB98106BDAE7F039D402E5DBD2CB8ADC5CF24828A100F602EAFA21557139D97086941F21BC78F48732E730CC8813B06C3F443E8620BBD5A26EEFA324AC15D41BFBE1540A643C2CC4730B8D77997C1D8142EAF99637535198EBDDFD2C8755D402BF97D39C6C194F22BF9852AA22D96E2300C9D49B67895DBDA33F59B88B5180A3A95AEF36F2EF2BC03DC9767E32370772464C1E44D0BABB4F67B6DB51F718365F86D67772A2BA4F0054A4CFD24A9EC81F459F6605F3E7EEE3C3953BB8FBFE05D5004B40969DD6A6008A6FE40B53CCDC8A2FF5AA977F106A7962DE2F8563277EC63D2FD457B5EDB35EE6E081DEC60A98DF886B99A15E2C23127BBEB4F01F89333440ACBFB7E2C55D01086A325C665DE8B9EDAE7730049E7B4361B21ABB1ABB8E81791EC82DCE3F1DDF0CFB626020A61D603D125B64E338372F5D0A64CECC4F456AAD3945B84E295DF8BD918F932027249D1012BFD4E65E4EDD444F55F4ADE8783D70D58CDE8FD8693E3AFE130D0834FD291AA62272FA04AFBC3F83C24444BDA85AAD864ADA7CE013E402BDEAE481435C448E25568607D2D4E38602C5551045D42885709BDA53C15D11DBBB3064E8290846EC59DF48E82324AB65D378A92FF93CC21BE4F305D6D4F44AB7CFA33FD97C457A70068402154059910E04031A284837C4BB5162A046EA579FB4D0B84BB88F8BC0762D39E877A8E86CEDE90A7E135CB80A4BEFCF4E4B26F77C8698F7F4F885C2F95B5171FC59FD844B12169736C62F89928E1FFB5F400E0B8D6DC435EA26738A076A68F24FE792E5FB8AA811EE75B7D89D5C6CCB2FC2B3C4AE2050C2709DFB63D308BEF8A2811138DF6108393C955227C6E928511C36491585B223017633D5B4AA52F69021BCEDAFB5BC8D966371D5C90B597E4083EA0D31FA856F2AF8AF57A4639CDC8C336572E2AB89224DC8E2B03675B6A7F0E9B7737BE944D69D908761841A1D8FC9B19E7B57D27AF514997C1DF39EEC0AE6A70E163DE86C242473D75CBEEEE9FE509FF4A52438402E853EEE7C67898641A86F4DD834786E93DD06E0555FB7BF4B305C19FE3654D94DC35642B048F590F2BB7003F3093C29F30EB61F5C0D894307D6E22E7593903950184C2188E4679FBE27759DD76C2783C6A7C19F341E846AF95A657BCD30F633F0200D78A691289CD5C4798B99C30185AB7B0212695C6D4DCED173E475FCCE7D287B0D620A16626E18BAC9BA0CCF289D229C39AAE066B436655ABCB333DEDD3FD751F1720B88AD36422310E8E5B0298F8D1A6C4710EABFFDE6185CC222EB02542013B369417CED1A318AF650F1D651534490D90DA00727A8F0E360C05AE27129666FA3D2D0703C3A5549F5F7F74440CAAF3909B2282D6B2941A831D32C95B7DA54507DBC134DF88599C67A5B0A9D13236A68F35E37BFCD54C113BFCEAF88BE1D435C1D49D03704494137197F1A7220B60256C7FBA1AD5B5868153743AB59E2E992C2B77AC5924781ED0CBE9601E6D6EDBBB4BAD9C91FC86722E9284BC0D232206E67CF45262A60110CF0E70494F55059EFC5D8024A34FEBD6C67A1358E168ECFD8280385B241045EE3E7528E883E69549271D715614CEAD273B71E87F1B08EFE8A2D8BD36929E13DB3F7275BDCEC1C4723DF334B4C6D91450D6A62E7B707D2390DC1FC3CA110B7B784833F01AAC28947C97B90871FDC0A150D44EDC8A62B4C5ED42A059CEEADCCBB8C32F44846DD3A96FE7D368A60265BA3722A7531C0ABC7FD0F0E85960374E29CA36A4A12F239AEEF40DB0ABE093DF4ED08FD03D5958CC70D8186FF2DD16C336850B78C1081D4C507D32D4F05D290F8385689629E180DA6507B2D34FF30D445C85814EE94119B9BF66242850F2A4D5BB3CD025BD75A21433DEE9C27F4151FEB309574C9DCD84486E2D21AE7881CB4EAD4CC5BC8539DCCD0094EFF373813EB37FBAE8F0EE83B8A7E8AF9C4E24A11115CE50D9227C2AE83F59800BD06809AE120B5D75042D1952572A9485179F9A76AD305D14E2BCA2494835F1492E28BA5DC58F86AD401EE7A737DEC12CF92430066D636E23E273DD5E8365F7DE82877A71F7465BD9B367F644C2DF0F869B869A265AC716A36C8A79C0B5F4F760DA09F4892F5A26EA313642E1641FBCD6EAF4CE96BA124C05D6B02EA3ECE8CEEBBB4B5ED97899397725DE7C1BDB4FA149AE1CB85048E23A09958236E22034795F028DDB21AC0C08CF965D1E2DF91DC2FEFB003C9AA9B39ED1867C6A761163EAA9B3DA584A44E8EF78D1771DCDA4E1BC70E704452D5AF86F01E417A5C8D73680CC7224300BC0655CE88CA33D3FB01BA51C0DBEE5B10B8FBF9B903026AAB67AAF96FB4E08424DE13F355E5891B7C0D7AE1724AC1B7F13347B9B241D3B6E578442DAE06874099BB50B644F31CC9B392D208BC1D3280A7B6A6D734763B058B65874EB793EF9021CF449621803217FAA47A8047E09AE197474E030C04C29D508876C5EAEC6E8F861546848675F04321A50EEA22A5FA392121C55E52C59352425D0DACE589AE75690B8209301ADF3B00BD713A17CC1DAA25A65E4CC3F7DF32140D31DCF9ABA0168971E20A3B13648C345D437023C16846A3EF92E8B75451B2D64C27B2631100C816CB65141E0F4B340F0826EBE11DEC77B66FE209C27E94BBD73B4AA02B303818D4DB9E7C6B86F33753FF9563C7231342EEE362BF662B21CD64694069570F0A2D7F7B7885A3C777E4128E512C69824241B7F26DA2FB4B92512AADC3945A720773915885E4AAA1F431CD154F1C883E419974003A3636F4FC84121A7FB87C208495449793781C7D524BA44604D325E6ABA53B05B6E0E3ACC6EEA2E28527DD65FB30F84981D2380FEEE1CC50A5F58A76EE76016649181DB08E363322E605406B825D8151C9A85A02EF9E07FE129D0496F23A80BE450792AA8AF299E3052FA63FE5F6BA576B0A8AB5187C33589DB38E5804882A02CEA61E88532620F64079748E54878B6C15C72749FB9AFACF876A4EBC79A95EAA6B0C03A6A9BBE781953B440B7AE2EB030E2944568419954D2DC193E2A274D628026261B8E4ADF0EC20DEFFACD1A9A3B8380B01A2EF7A2241FE4C26DA3F4FB41A29FFDA50010423E1CC3EFE7A17D5F0BE70870CC4D4CF9CDAEFA05469EDFFC4C9D096B4653623D6939E0AB1EC2A4CD2EE12824EFA25FA665921A1FE97FD7D445A66BA929A94F1013DEB6C6B008AB1F5D8DC76E4A0D87A74293DA2F4EC0814D6F686EB71D6A65E432EE20A7FD368A1363CEC6B3171ABF0B2E91AC019D9455ECFCFFC50B887124316D9425C9C241C3A91C356013FA852F4A7D74265696D1D2CB1D7002283C2F2BC435B8514109D361ED63ABDD26C928D67CE29BFDBA0F166BEF1B20A8A329E78CAD19EB2B8D13C4F58AE0DD26BFA7B18850012E485B89A54312C91EA862659209DDBBB287DF1864AD6F0569E774F4560B7A1B2BEC969CC841825BDBCD357E6C16A75045C9D54DBD0021E41D47A09CCF70E9DB766E5A981D402C28A183D06F65E8F4A102D02E9EE184162DE14C5D5E6AA375FC5D62244C42358B9C6A0F354A3B1AE4F00222D43A38EDECEA52904A264C2694A43BA86CC01D80E295107DF95CC1E82AEE5049D764D1DD4AA1C0631D175843A678B4A39893E24D0AD6FBA3A99FCDBCB87A5D3716E0AB10AD03589FBF55E02B502519281DFF9D14BF0B71B713D98F620EF13536F18ED628F3A25D206325BACEA3D4FFF181BA97375F39410687537D159B2CBFB8CDCA44CEF9D0AA9921FF5C0F59EDEF19105B5117EFA493BF651165275371E5929F4048B9CA52E2A1F1EF95943A6812B297F5E9B8727CBE15FDA87EAD75EF607C310D284E63721F8ECE0292F23332CDFC02642595FA9A72C448AACCEF95B0703B3C61203B79150F9688FD81CADAB3355160799CF1431C3526A82E48BCA885AF4D4F1C7BA3573952D11C6C63B054602116600D3C30F45FE90A352033EA71D87A81D1684E5A29DEF70C6F72AE5A004D3E3836FFA75D7A17781E10F73A4FCC223C4F2411F6BDF6AB46848FC944ECFD0419C8BC389C084DBCB7CA071B1F87D15BA3FB8B07DE4537C7FB1B1904D6610D9EB9C64604F2373580CC7884BACE6D3B48A34E043CF0A612E9ED9C31881FAAC71940B6E034992B323BFE1799D5CD5AE8466D79DE93F50C457F44BC194A7E89601D9836FD723FD2899D22D59A9F70B83BF0AD8D672192F9E97EB36D7682674124CD2F3FBC71DF5BA608088F4473BD8AC49125D74EDF57CD1F041462704195A0F049E49D1117B90681CDC6C968097C76B8E0E9B7D280D1153B3E7C88AC379368690CA4B44DC11EA323961182C1A4FA1DA169D1FCD55493B937631F1B71A820CBC0F05158620C2C3A46FFBC536D5EC093E0EAAA690687530B4C59429E9E5B42310AA46497A87A0043B7148408433232FF31D722EE34455294FE647AC02D4222F296244254188219741787CFC26E744CCF89021F1C0A9B1C9418F04045B9555B569A262D444188D5FFA0F880FE1F14897E4E5E4E3C632ED7B30E77F2A269BF9E5BD028B4ACFEFB46FD06FDAB197CB38F8FB6E3490CED668077C6E4FDE169787F640737448952C862349808390CA81946B0CF1907FC9DD49F8A926CC5D5494AE13B35F27D60FB89167E41DE5F14DB5306D02F8A13032BB92712E51B93E5EF55865A00AB92726CB848D00ECD10B5BCC9F84F27223E9B821F9CD8E2B34EEE572071025B83E4E492E4915CD6EF52604D0305616CBFD3AB539817B6E939E5C11D33AAAB30DBBD6FC0FCC459EF4CD748664F188851F62FC123AFB80AF20F5F3D2D88A2B324DEFB8ED89E62D8B0EAF2FBBA8862A713BFC5F0DCCECD86F366FB1F54827890C301B5C67422842D86BD95A158FF2E4851B70F051795588E1D167E796EECB490B13E417A42AD1386C0FB88ADAE96EBE8E6D0C457A76B6363E9F301264D911FA76564F14E9D83307D191EFAA488D90EC0B5F8DB1763CF84353292E32D3FA9CF296C3A50721A94B4F4196A6E7577E28753C5DD31963101D8E1E91F72CC666A7ADB525B465A96106F9653A499170D7CE80E414C74E9C47601AF53AF5E14F47CDD099615B6D6D8F7068B5B902A3F2E72CD79CC177E1ACD0306C3D3D517DF3D0CC83998478BEEBFEF42C09C7C8E2A428F509BCEAB30FE3E030EEBCE1676BB0F549CECB2F2D42211991EFDD6F3BEB1F9EE148162B494E44BBAC301660055F82FFC3D6CDE5A15BC91957D7C91DBF99C42F801AB64223ACE4EA0EAFFAA74B4D215080180B18B0D921D4633B6703C3689C9D9759225F02949E48F5E3D4557BE3FD4F60E47A879497A136D732F96A0A33D5F75A1497A1917906EC7B2A5134680809EE9D0F544809F5BA9C7F929F0217C19D5B33EB7EFF98D218172989613C1D521E7FA64EAB4AA19DAD0BEBAA4D7262DE2081A9DCC0684D3FD32151B29A8124435D8AD22D90B4C0B754CBA2B239C100EE68704D1F94C73E8CAAC0BFBF4C079C113D0DC310C25CD91495B437DF82AE6A892F13E04413B70B7EA4D440DB6A369A1337E14C0B8BCDDCE92EB892161F355BD1E656D2E666F8C07E62D3E9F1488B9F8C746399A28D981DCC4F90F690122DD0CC395B9E2CE9112B9A130BBCB72A8AD513E3BBC2F0E5F86F8E91D490DA05C08F20DEAEEDEAE9210D7DB339A1BF7B990F8CF0A35DDF0D55F2AE4D600DCC53F7B517C7D29C05C53874839949A81DCAA7236B5345504EC481ACB8B6A530CB29997CD086F69E0DEE4F731F354C2C388A14B96155F94212FA04E9C40C3F899A3E0395C15570D05CFD069B7DF13C524C75D692DB418E773CC3AC245A4762D89D930EB92EDF3D92E805AB08F7F1EC73D51666959F1450CEE5EECE771D5090DC6AFEC23F40B3B14E4E1EBC5B0AC37EC79593C11541799DDCDCC8442A6213AD1C4B64C4C3668A6D88CB0FFB6B25CC0F192D3DCDABF3C6D0D358FF2BD223DDAD52E430892C46E49500F0237AF01878C5E2CF8B5416028D093F12F2F5DDD9CBD395FD2F141B24CAABE9DDBBCD825AE8050724CBC344F96D8C56C24549B0F46D5FCD16375C6BA7D7AB366CD9C6A00136B87C56C9C62A96C8F5ACCFE742ADEF467701D882464051631FE2223FF6F95BAE7A5D1C4D8DE1DFD8E5A062B18C3BDD9212D922B2B20BBC06EF3F932B57A568ECBCC6082A46182CE31163B599EF5D9A150BD505B50BA09D9C1CD310001954F6562623363BB27CB48ADFDFB2F71CBE6DE0CB209FA071B9D9E111A03263B893704B2299155B010A8351FD4039217BB55555D58E09FABB99C4DB2351F3225D8AD4D514606F3B85B398A3D250DFCF66A129FF65EB08719105A74E25100C8E07245E5012445F9A762F6957835E408B253B440C4F6A0F89BFD300B3F52BC2CE813B131535C59D6253177EFBE89CA8178432FFA18F2ACB9F1A88B01DA73A72A206DED6FF2BBA630F333BC453AD328889A671946FF03BE23DDDEAF343EA80CB033A8B68B3C17135D8AE0D21548BD77D675BFF09532A882A3E44D88F17B5E698235606E9D8A55E4A597A2E195AE6372396D0FA5BBCA93132A2C0806DEC625B37FD2DE028449D7F5A0EBC6FF1A1E7DB33997E7FE2365D46AE7229022CE491EB38AB791B45C8BE9B6EB1BBB50906C4D2175EE829A36E515AA07F792538A34D127C931153B1D6D859D34593DC25149E9164FFE81D58F6504E2AD8D19B8EBA0DCBA5B2CF12C5F11C9D6AE06B83D6C1C1CA5C9CF8BA0E0A8D11EF7CB6854F902B98B17D68EDF3DFA2F8B7499FDCC73D8D6E71AFEE17562A9CCF4DC761F11EFA8520D13112F6B463D88849D5316ACE61D3D764AAB9ABD5066533D366BDACC9FCE60F163842129EFD7C7F2685F67586FF6AC9711AFE514EECFF2A722C3B38D2A51C0BFA90D7D575708938A2E86F77D7CE9B729B19A6727E4E9E10D4EBFA81525645F6DFEE6A8A05D36867A81798EF4706EA2C4C8ADC91D5969EC369966972ED755502A8A8E648A02A1DDF0B07B8AAB31CC15EC2E210689AD307D8AB4B95356DB458FCFF5703C164D71BC4C9D0186579A62517E35DFDD88712DD8520F03FD45215E2C9896CB19BEAF66323891AC379C13F246BE05EDA623691C071D66EFE99864F9C94B33F1D185D411CC0635E18B83CD8E167105D64923F7008094F8AF4F70D4AE88A832BEBEE3B57C0A8A1D45126AA73C9AF52D2198CA39556F23A01C218F5C4DA8419CCA11C1BC689A93E2390440752E579F177AB739E1258AAA48B60A9A2516E82C517CCF9AB5913F82447096C6E218FBA8929E4C74F3B637DC7FB0914E8F506A410EA1DF12E2E674FF0CF6A9AF459BBF6B164197AE87355C56EE1DA41C96072621716327DB9B4A6715FC7644FD43B0B70735EE90B7878F77C7A74630A366366C990E598E9A3DD39ECCF8324504DA49FA54A3EE7FA0A2B90DB9DD7BD3A29480C13D1BC230740BF6F9C50C2CFEEFA62D843B0AB9CF1CA4415395B1A94F0B73E2ADA5B9B21BECD58529A2919EDE578C36CE1247912C88436156F57AE092A9ED06A5462497EBA5A5833EA46A88B0021DE82DB190D4EEBC54ED5ABD13BD2A555BD5F5EF3CA0CAE9E323B2F7627986147FA9ABF8B289895E93D8A7B0B8A5240F0B661BEDDA10702DB939B903192D75A709692784949626C41F2F4E8C79153EE859310B32B1EE8D1F5CB749DFC1523D4EFDE80A6F2B0C677247E3635BF629179F2F5AE83763B5A3EA96208504E937DE733177F404BD83824D85C2E149CDF280F67F180B381FFE02EBF9AF08D4EE7265F7DCBF0CC443C1FB054905F2CDE5F37BC09C0F9BF28F84AAECFDBAB856F9897B1C33713EDBFAC4A296C203ED2C4E427F49197276D1FE0DD62CDD36022B7BDFDDD3823D41D856694556199EEC522D300C848A384E37086C045876DF34CA54005AAC7363903F2EE222398B6507823809D9E5DABCFAA0BC74E1D133368AE5ABA808E23858371C81A2DDC6AA8246D14421F489B3D348BE0C3F348CED185ECCF972FF190CD9DAB3FA2754DA937EDE81BB1DB6B5457F382814952AFAB4907A7BFF078636AB275873612C83630A1D1D42332309F58575662649D1A17D7B51FB26BD40E514377D49584344E94C4F0E848339F6356ADF7B42D7E320CACAC72F24AE67AC63B23864CEA8C84F6DE5754EFD68A0B1F24493D2CB8AE10E0082E9AF35032475E03AFDE1D818AD7E56CA741AC13CC5DE4C4DD0575AB8A0BFAECD85951486B28DB5059B4E53BB74C94C2E09B50B270177376064A7F0A230F87D3D2A55FA6979035DDAC3F121A7F91E29DFB70117A139FCFA936182D76448079914EA3659E65009848B99C207B0F1E3353CE8271AFDE1FA38913AB5EEDD2EF423A3E5103B6FB3A00972F0D1BDF3EC415E6DE807EC7D59A9C255A581F1F90CF5D8A86D5D569B72F348A1BDEDFCEDECACCA52DE88EFF8ADC5841EBA28F156B5E7B5BD68D154B45C5D0C9F065909FE40C0EB3255A4495DAD3D75B7952C8115490A742BF546B20BBE076710D321AE4527DFC0C37EBEC238CB5335485D3CFFCF1E808D68047D1810BE4E122C63699940A46C5E92DB9B030FF6229CA7613E6C37822CEDC5B337DC44696F143CFDF95FDFC078B64C505CCB20F3819C5FFD63DBD46929F628AEC084C0DE542EF0EAD8A2A3D7935BBF370DC75C2748BDB6A59A107BD3BAE84398DB88C7458A0FD5DE3DA574458ECD49C7117EBCC54A84C2190A3D395EFE4D34F3100582EBCF1C88EACBC526E3AEC1A8E75208BE452D2691D028D80D02FC1BF4C6EC36647C56FC5CAB7F2D48249E2738484DB9FF17AEC4494901C625E76B1797006C642F63A34B22A7730F368AA899CC7D8A142E60D4DE75E67BC872D8E83F5666CC8321A25E3542A0F70D1158D0F5DA76C4D8CA08B13BBF1B09216B0A81714B4860E46857E351C7C99A43ED162C7FA7E016880B5C063BA00DEB64B793F5BBEA439297DCCEA01AC891BE5DD2BEB3F876651EC868FF0163BE6F1E8A838E6B7C3AA63E2E4DC4C49DD48F53F913002D6A610474A47E1E39764A928D5435A04B9A60D72416368FEB41308569342679E546EC0F60D9D81547981AA4A8E4E7E96A56501305B8348C26E187BD0979D7090A2E3F893E2870EB88390F14DA2A00153C2CCBB309D38EBBB2359B9317F9DB1665593B023772326814CFD6F589DB133377D86B2CB05C869A49052FD2DAB1457FA7FCD0EF3DD3A5AC7147AE1838BBD109EB0CDACCD9AFC8A3AF15794F54364F82FF25EA2346A363C4DCC73DF64E6D88E36F919A740C1C4CB7C8A3FA50D63313D614815011F14F2115EBCAC93E6AEE230ED996B7AEB7194AA05A5E951C7C470F83C610A3391F2D609A0F667D41BB67E99F9DEF0146BCFAA483FE337CA284582AA3BBEACB761110DD048C52B2D02DC7C4E4183B5D3B469ADB91F14B5EB5B88A42977613E50336309BC00273561150DF9DFB3573DA4BCD65AA2468293E4F8428A4B653D8230A230E199071F968FFDE1F47EBA36DEDD5C228D98E76D88C2478774B057CFDCE32EF80CBD96C142976048B977C900C7C8E228AB1AEBF885D68114BFB760D95EB4EA115F78484B746042CCB7407D891E94B52E04F6C1A3352C39EF82B2FA2614DB946A2A916B44B09B8E4A02EBB7F0DA4FEF1616C669F6A66C726789C32550E8D08B55AFDC60A18786BB1BAD215E7DD6EE9AD421448C0226809B40900E4F8ACCF756603B671BD5793558FC036637CFA230D725C7AF1148D5B15EA3E629B1544EBE18A7FB90F14EDC8EF20619CF07C972CCF8CEA8ECDF63A78CA374C47CB4C7D2B88DA2C8D60C3DC3568DC969D8E788766A9E7056DC09B891884FC1081C8F7E320384B26284EBC5BA09C49C8C062304E9C81E044A9E30410C921AD56DE41D6CA0C8DDACCD8C4015B584663562F5F762FCFD88A9883655FAFEDD57C830A4C12E75CC5F01616CFBFD3E2BE13D9849858F65BED20F7740031BF456317BC6FB84B95A72A072022F893BBDD7DBF7178AE5BC74B809E584FB9F8370C271DE71A715DD3AC86E9D49B7E1DB31365BDE35F4381C6E92813A5968C04B2BA82CA33BCBFAF4A434EACCA17CBD30589C31D5B9B1318DA9E1FD87F3836E03636861A538CD133B2E4282703847CE00F2C98718B58827321655FF29D7871F20EA5432EDD7694BCF66030E69DEE2998A067EED34A95EEC1E70AD8E18906890E70B2E65035C003C5F203309B392756B2CB53AEF6B21AFCBA320E1053678ACE6C9D93CEEAEFA99C3D0FFCAA9F32CBF7F60A3F731B0E7F98DBF15D301AFC2F69ECE102CDE5E716A98766C0F82592EEC7A29338D0A146E2CFA2FF2505DBDD2A9CBE3F30F00DED8780479CD4CDBCDCA17A6497514363115B63D67C960E4CBACC525291F55B5FBA30C4A124AD47AA134AA6BB27EF1A55E77873A6F4716E46F89BB3F9B159D1F1E80501AD3A967D4B57C7E390933A0CEA93E1FB5A69DE53FAE3541D974899F276BCA239C4AE553940EC02BC56C7B5B9628F384E49F02D1F12D0C67B554B0BD645A33459733A41B1E01E73429A45F0B47AE9D1F1A92D487D59322BC2309396867DD65A96675958DF308D99D9FFA90A1DD78FE382E15510DDF9E7B92EC732FFDBF316083B4EFE3C9803AE2DE9FB15526A6D023C337C5ED603C7A242D7A995FAC76B47FD4D07CE7AFBB82489CDBE44AE886DB161904BDE73670DBCFC26276BADFB156A3AA69F9E69A52C7F52EB88FDADF9F3FCF5567252CE550572F1E826FB29645C173DE642517EECE17FD8AC02A68D143023EFC0A9D9F53644D22933637F5B2369E6E32C54707AB577D2990505DCD8D871485B9EDBF58A44FF84413CA20B711C1AFD8586839445585420573FE627EA14D607CE06F7E505DE6B5E59D4EE988CDA3ECEB5862D8C5E529AEEB3CFA529722433600D95DFB92217DA598395EC4D525F4109C5C91F5511B999263CFAB014C5B716B443ABECB7BEA78D6B84ECE3A43850B08BF194449BEE2D0432D7D938447ECF784010F1F5A24199CB49507C1D5A2C7B4FABDAF39B41B3162EC6B38AEFD833A30C488778F30204959F05537BB516AE4B4D259B3E5A47305482ECBA84F4E6A18230DE2320904B321D32DE58626D4B74068959C1390B043CA8245AE6DFC04C70F4BFE2133DF0D00BBDE3DE363EEED5E6C90C78018471CBE2C193F5C5F9334AA19FB11C6E096330117BC074E708D7EC70E40B1421C255D8757E6C795C804ACCA18C115B4158F27C6FB3ACB3E6981B25A3A3992B0FD90C8B49D39157AA18A79CBB0CC934835B6FFB678C3F8B1871C655B844689DBA1040CA823D8351997983C17B0532A50CAD2E92438502A8514E16793E32246A19A248E4D20FDFEAF1BE386F92B79440B87379650A33731A81101B22B410123292327881FAB6AE7C7FAD15E21D326874BFCCCDAC44499B8DA9D1F45CBEDDC47A2D98AF6C4A0FDDC76CCEE140740C9FE0ED7E8D5A3C523DD25D097E3ED991EF1D1E74B6EE71B52006E8DAB83E971B84E865989FCF98B3B7F142D5DE6D9BA6C4A8B785870ED6282C9BA1D92A8DDEB22F97C4F3A4088C6D0AE523D41C676CBC8326CDB8ACA29FBBD68803BEBF0A78C619CD392A65824E3D550F67BC13DC15244D81D1107E938C60AE615A4C4E699AAC053CB57E5CE0ADDFEA90D17EA3450DD9B367ADD7B77ABA87A30808A51C79DDFA5D944778E782C640685F4880FC0CF22B239970FC00E33230AA5B2DAD05062699CD7D1BCF3CF3322BB2DCB357E441C5E5D659E3F30D3A57F9A1C80DA1588B4A60DB821A3C36EB89D621E870522A325ABF4CBF345823211BB2950ED71F099307119A144EDC77E98B0B9DF69C398BA920879B7EC82AA03A5CB1BE3A9E6B72CCBD20F6902EEAF7DC69C6E5A9D3C3E9C25ABC09F0F232F15C4FB8A266232460416D209A2CB105825B471A22A2E806584730C85BB255B700DCE37B6241453912DD69171E1B5ECDD70BB6028B58F567C77F74D391748150240C53B1955927F07A5785222C7C041C1C1B7317630FEFDE8C5C8EB26B0358BBD48AB3C585D7552DE85512419450B049D24C3009161A2962E08FB916C448202987C10F849E7BF67B295FE2249D67577C8529FD602F463566F7C488F7D81E5E32E7E85FA85F728770526A4BB922E99944EBD07B7768B425D863EAA799BFE49523FED35E1B4BAD9A81F26D618D4943069339D8EA75B1783AE7B4B0E3EC858E9701CA29DC8A7F22EBF3F6207F87B37D3B4AE1792D780045F3F57CCE6BD84A14DD7D2D9B5393BC4D74103676C18D7AA8BA08BF03634B56947C2D7D34827F0E69EE32AAB27C7E4EC57F7765D89E56951FFC03C8F3DEF343A230240454633806A26E4EF9AA56C813816A139EBCD6FC05C3531CC45FD9D2F00F4894DDC5FB1D26EDF5736674CBC5FB1D5CC0343B20D8C85E042CBA37F9E571BA6F614C04D65A3F94B5C85B51E9A7CC742B9F311F23458771716CAEEA6BFA1528BC02B44047F521650985922D4AD1FA55016AAD8B7034B6F73316DE91BB80BC803488FFD367F5676C9C9975B3DC61D0523B126D0848F5853F7FBB85FC6F207D045EC011D87C64663AE47CD9D0E6A4DA5CD828CBF87A8C132889412E63DEFD2F36D6302D24063B972E89BA77171989054441BDCBCFC8A8C12F9ED7719F97F8299F791493449BD7A5A0F0288E6EFCDE91F4E2B1B1A150CBD71AF2FF34ADBAB77687B5AC6C24755F696790F4C72006AE10D203754366EA6E4049D502B1BE5BABA41084BB298913FE4FE03A385A440C3DCDB6311C947BE102520C9175C1DF5EE41C49B4C7CAF913DB16E35BB8F0B74388B22364AF9BEE986F065A3B6FFB4BE446559744A2854670550868161DF4F6EAA7F57D8EEBDF34827DA13687D3EC725D62F35865F8BFC6B0260B083382D85BB6CB87B87E2FD38DE6ED1FBEBBD97F10F297922335A2B1520AB35BFA2946DEEAF2C117A0F4C8B395AAB717AC359FCE6BBDF39C8E914F5312A4993CE173F204FB72867C9505CEA27000BEE64ABB07CA04AD07C932C391E7DC459F8416A96A308D07F70C48AAB46F5DD14CBDD12BEC38E571C0273343E9E0E0FE19CB7734F9FB3E358E0A1DF1247435DFDEFFD5CE4AAF25BDD72FD8404CBC3BA7BD4E13BE224BDF826896293BC799E9ABBE933C3C6132E6AE412782720A74DFB219CFD4D764DB627CF2F848DA7970D4F0089B2C0B7565F77D3D279139FB9726039646DCED9E332D8E85C40C83BCE4372592A2AE641C16EE9FB28DAD7A5B77BFE468A5D2A858866A753DF482F39D847F8F50BF62B880CB3202D4BB4430ECCD526DA0FE39F52D8D2B24258FC666984B50629924FD97A6B741F1D026315EC953B8E859D2CA643975E7A795FC90DD5E96903ACC31F18BE901E485A01722DDFE51420FE5A8C4B7B472C9B9A951A557C3438B1AEE141B2F38DDE550836761451285FF6CDF80F5F823B55F6B39722264A861D9A2CBE08DCB9891791761AF2EBD807EC8A6EF9782142C95DBB2953099EA5D852524F6D3B9D388AFFD2E98B2228AF6448A0BFEAD7DB2E6EE7FD8B0D42B24D28358245537C717BBF4707CBD1536293C5940E236D1DAB210EE04C80845E75730A0EB14D3E1EF65B4A3203372B151DD98574D8E647372A7E108C7F0188CAD31312B6E784D68652C49DD912B07182D69D28D2146501F7968AF51320AAC0B77A1504E70536B3C72B6913B35B0E3F29FAF5423D9CF51B0EA71D9B16397840EC5F7617D4C0E204DCD58BC65F5CFB6A2FCDF71ED4F0297F66C21E4A370FC821E1373696EE085C43B6A138A8791F2E3FE080661AEBEA7D92368754682ABFE5C3E5CAE588D5FDFC80C2D4BFB032D28FAFD5F38418E27D1E62E98DED09E6D6E5652BB4CADC4EED8DFBBA68B171901474CE8F41CBB399973637A5240598CDF192C7C560E60F4B4D289C54C3827A23AC49483D5C6BC4BC1861B0E54483DC12C9334F2F5C0B0F18DCD3F8657D129DBA05A8C161AE2A64CB5DC70292C15449A37F1C227DB40F882AB0EE1C128FF9306010DDBDAC96AB6435FFEE070ABE036531A8BB4C7E244BB1F8721B4AA318C5A2CBE53B207870C4340FC9C10D076E42AA77A4D8D1E360AA461EC0C8960726DC1B9169CD2E9E14710C0CDEED334FE2F781D6655AA140DA2B3ED345D2A482DCE127A9425D445D61CD56A152A2AFADE3A8A2CEB63E763E9904BF67F521968CD892FCD221582B6320A30DDB6BBFA61321FE44DE8D5012938067155E055BAB018ACA4DEB79DCC2301F1970C572EE0C4FD9E75D14632520584017CE2B61F4581CE186135FA5472FB37381ADA7E93CC712D0C725E437C5514A5AD3F7A60CCF8F33CDAAAB9569A00983999385CC46CA26ADBF635E6135F0559753DEBE4361FABE4455A9AFD64BE87E41CE372AA6D013A51C99FFB62949401CEC58679E70DC27261A642112532AFD8FAB14E9D29A18066166834A88AF360E0500D626B9166A0BAAE65DC24BB32D901CD9EA04D8712976809C4AA13CB69A73F33732418E7645E34CB690EA875D53C06F4F6B7E5AF4FD07EC629F72B6525EE2007E8D365BB9B7992B937C3143982B170F93F439443153945B0F6350EB3E49F7E9CBD3CAFE17D5F0F5804F7B0D2FFF764BBA06EC3C10828654FA65A7AF4FA3EF2D42890E6FAD9D7AEE5F5B9907EE50542C3356ADB9FF4637415BA6F9FD72289C6D4692DD18550008E5D22B307664B6ECEDAB92875F3C3D6C057BDE57299D7E035BD2C24ABF46A4619589E6B0FDE1904C784F11A9AA652CBA06399DBD66DCFD08F98E955F081098C2D1DB0842C607426C06E4565AFD20E3FBCDF3403D195300693B98A4F074A1997CF2CE95D0589A5DDDE5AEEF8D96EDFCF06AAB1C1304CE0D6F9C2B3F18BD3B3936A77F54821013088008B249827074B86E8A86BA446572A64D9D79FB8B772CB0FD00C0FC55F88989FAA0978A3C4CEF406E6F361A0BECDD1551B49A3F8D614668B174FADE0C85EEAAC5DADEA7642CF0EF6E7A37714F7D782F3E0DC81F9F238A9ED75AFF1F86DA678868244E7078AE09EE5A25432DA8F0FB47AED394D83B2D0164CC7EE2400AC0E2210C41FFC493C7E9439760C2E928F2EB4C89BFEB4FDB0E2CD7D95B797F84322372E560F707ECFCD4F08FC75E53063FBC186AA1F1AF0DC30DE3DCFC5CB94C6C6891B9ED605480A10ACCC9FA4097C56B0EA5EFF360073CA4FB0A8122629A5D98F1DB53EE140FCA6EF7EFDD6B041C5D1DAB6CFFE9465EA30E481EFF2B2902E8C11AE08EF7ECCB51D69626D7601C986853F9C191CD33E796D68D3E272AB9F9D47A93A96C22281F7F6104A48954ECC85C447A2FEE8D20E04269CB0CDBE8F8182E323DF40D4386318D7071CA86BFFF2342890B51CF637A75BDA2C933246FD0AC10C9EB4F81D15A8E1341864BBFD69D5F0E2F86B1DAA562ABE6094B21A5CEDE57DB9E0424671C17897F7F2B978E6F497DB924BC8098CB191FE9B6067E5B6EB44EE51FC4C2BB6D7A099F90424769BC1A5E5EA14075BEC4475F46888FBCCB1BC4BC1CD2A89A9E065DBE15DF7FC9BEBD5DB234C59B3282682DEFDB063976154DEF92B386C89EE76F22D657E11F56B4D23172F4F84BB8A4087282541820134653D2CE2A53629390823CD5849A324A3949B5E22A534BB582AE7A89940E0395CBB40AD3C9FCE544631F1AD3F42023936B8B4C940D36948B132F0569D84121093A9EB27C59175B44C5AF37CBCDE21696D698C3B14E723C686253E0106FD38BE4AF40614F08D597FFCD121EEC03E6E082EB8111F1CE405AB16542FFA0BB707A42CEE15670C24F39B3BF653F08FBBC852531CE0ED9E1B61A242AA6B0BA17A6EE163C8A8650F681607CEDF7784F6E1459DBEAA9D7D5B7BC8AFACD5ED4C9F8945FB136C3127E423E3A8FE571BF4D8F468452ACEA24239616BA2BF12C4AE9CED0A1A7262B4FC5F26E709EA8E86E83BDD1763D4BB4861624108E1B031F852F2016B530F71F7374AFF33BE561EA29414466645487D07F52A8252EBA0C7D127E253806D3986B072655EBC49E3DB5D164FE723B1F88BD03CD12FCBD9422ACD3455D7EDB36942AEA2787CC104F77EA390390B664C258B8B8F158DDBFC86E04A59E63707B62F4D375A77A3389DCC849EFD31D9469F84232CDFC92C27DB95A8042B7307B0D2C8BDDFDC7205F352D312AE1C6B43928400B5328C0CFA3E5C0DE361A208888DBFCBA65F396E01FC26014E15A37EFD983F2C3F84341FB94E5D4942A1AEAFD37061FDB6D48BDD33BB0441EA03D7E6B7CB315B9305C73475B76C8AD188973D91204633E3829A776E4C8041E199E1B90C73305E845B2B6CE1BF004ADE37D2D80AD7D81BA172E7E759A9D58D6F80E1E3B0932C80E8C6D841FE4CAF403DE4E94F4808360E88E6C01A44F832689B00F2AA5F63E45213E70BA3FFCEC6BD17F4BC127FB76E84BCCF74CA139AEF7CA27C41EBAE24C7E315CB722F84C8CDAAF0572F2AA83EE3374607B1787634722837B4773A58891BEB303A0EE0C1EFB6FEC4662F39951A8A6BB6BE397D4CB93DACD92050E05491129ADB10609775EF3BBDC1E5326F28CC6D183FF4C01FD7C2477D5DAD9EE7A379F2EA9B146420345F7E3203866FEB1F038A04324FA3E0C803F721A162835814BEDA94F250B63956B6D329354DE7149950FF56A6BC89A7AC556A4592EF34D752E515C676D4F47E0345107338D2DEB679FAAFADB33A1671858B81F245C963AECC780C4AA1F6B50B6425F7A6A132BBAA31193F4BEC3CEF96AFE37F952B1B8E9E9374443F270FCC81E6573481D973BF2D7D14879AC5020E672A53766F32194BF0C6ABB81E8C109F5833F80702ECFC819EB498FA1FE8B6C87942F0A131C8E76DA0672B0CB2BDDAE302E0DEDF61B5221F58168200C220A6EC33835C3A05EF5D4E193468BFE88F1F907383991D06E8E932E7C5869EB32F06AA64E3D35A780EBDAE91AEA17DF77819FFABECEC425CEEAF07D9ECBA42EC8BE375B152E8F76491AAC236F341049DFA5483E778DBAD53D9DB77893BAE36FDCE82A8017CB9D8FD9A8505CD260DD3E40D54EBDEC0CDF2A6CA2EDC2CB92404159C2ABDBAABF0E11DBE592C3812DE5F244AD5B367F46A52CEBE849BBD6C24EA54C8AF30CFF328DC918D0412B02455D6BE24C7E8A5C1D67680689692D8E9A282C49E568691DEEED4DE9E415B184DCD8A8DE9F74A85406DA571E45BFD8511F4C24BB17D26F4D4EEDCBEF02963CB6C96DD1060474A1CE9597E245216344EC9DC75DD8CFE66DDE51A00140550326C9C125252AD490D5529D783F02C8FD0B2AB0149DB8F4A95FE6E034997CD0B93C3949521CD21860105A4706F835647E1DE84890B14051BCFFF9BB20BA74234EA159431B3958599E1114906B107DB4F7767B8799A58F36EA3B0D06CA7A3314D1777B29709AE39F1744065E701A1B2C0718CFCF075466F43E531ED375DDA56CA0C42ED796EDC29DD90069B56CB8C345F55AA4675D47652A9107BD5F9DAAC6E2419540D04C13073618B0AA1D4EF9A48445E8B098D8F067C6B491A70B4F083E09A3BA2DD544DD28CCFB818EACB7E802A0ECDA35A0489EF272570D4DE8D7EA0AACB07ACAFD9493729BB8818E06ADC85FE52DA607EEB03F54FD6668AB514DFFABBC22E0B5FA85A6736F80ADA3EDDDA82AD0121922778FC83A6E62936AFC429F4B76F981EF7E9B1ABB1EED8E5901D50DDA74D9250F9B3DCDB493BDEE3D77CF4354D023D694058D3967F590A4C229C88C4F977C6DFBE844315403CB8A90F71EB8D7602BBBB9CD97D178695812DF4994309B5E3BACA663634CE3BC45741A18926D0AEBF931DF928A008CE7150BF1756AF5033A1F182F00E64827F272EF9A83A4E7DF01A4EFBB69EACD818EDF0E25385DCF858EF1BFD16696B77E3A1094B776D438E6DB5C8134DF7391B4F6E66F58C20B5E8F951A23EF8AAF4B84B7B2E3245142E6888E63A909DBBFE7C7C279533CB4C84C08613812FA86995102C6235FC505A50CA483F51DBF409C2AC07BA4E954A3925912A8316B8E0FE3E82656A62FE6F16E52138647B76CDC4871DCB3B4EA14118476D425C7778AE26D9D5669639622CB8B0EE21ECFA5485343C6D2CFAF65382C520DBA163596BDE88C8EFA1B340223124FD8AE9FFBB9DA87F8B38370267BB47E42D9CE6BB9C5D3B049E1C2656B59175C84FC072EF8334607C781F91925498625CED121D63C9AF44660EA19639169C8BDF61C7F31C79B9AF0C1BE2776FA30F3B4FCE2EC71F1D62EC8C809D1D4405175AE46906C963F8F5509C14B5D8E7DF93BF0CDE3C3DB54EB0871160CFFC18C6CAC6B7D1E9C4E68E552317FC60A9D194F3CE9BFB30AD9DDBFEAF87D58F72E68B10CBCC98165C5C85103DBCA7D9816210BBA5BB8AB8EF5CBA40E658921C534DDC653F50AD3A32CC2A8D70B779A3D8896AAD61068AF2F580828F93E8F6B5B7DA891452327C14CB12739D5773EE8D42825577F84A38AD6206E9158B75C471B7FB97C97D80C338AA2BB87B7C923897C6B83C9BC70C69BC77E43E5D0513F11ACF4AF4C84A20482371BF596EAA1DE24485701EB0F18FC1AAE6536DD81830019B49163CC4692D357D04249DE2B7AEFB09D8DCEFF295F2A8D19410817E045FFE9DF92600F8ECBDCE88BB3516CC9D8E4ABF23145CE83DB4B7AB67F6488E41839AC9AEF574A017CDA7B75EA78B4FAF9718EBD74A5E77E68D209F1FB7B1828ED61B4D1B9F7BCE7E1B7F0516D2970C8E3D8A96DBB0039DD2468872E5EAACE6A65AC736295996AE28EB0F10306CC421EB86C4F5678D84CA332C6375BF3EC854068E2B60BC636731425E4FEF6AB1A0F37CA1A2FC0EBC1B534FC7D94A430B174690126AF2404D353F490234077FF6603F49DF0B13EE0B2E13C67453046187AEB4857326BCD5BFDF8230DBF79A95177D28949F8F2FF47D0FE01AD0BF1D5374D4D753C5569C63D549C425380E282CD84D38D57B3B7F517F05A90404DB29A480058748BA13C10DCE68395D2E6DEF39B6AE1466F21C5993D8EED1583007657B6E0F5201B4677122FE1BF19AA14CF52A579006FFD84C718E702E083BFCC495221E76F706002F7A2DC599D71ABA1A0A843735BC415ED3DE513B240C46FC4E25A293AE850BB8E0A583B836B78ACF8EBC57E881AE16002B0A40236FA62C807BA346DA332A6E0D3C7FE563FB488AABF7A995629116A1F7928BE5C8049464CA755CE64350558538796CD53591F210729DA372BB4D0F5909EDF5D32C6FD73645CC840FF5190CD67065193388C9F2705003CFE6F6713ED8AD0555E059778DE646C0BD007858B7C39327F8E6C3B6CB0CC01777BDDC920BEEFB2E77743C9EDF7601A7D1DE948088869613994BD32CE03557FC4247B21754A919FD6C97C964780F1369072878459B8351ED7900773B7D9F710E7527CF399FEB75E3E2106E52C9BAD419441F0E2C7BDC05902A97F5F54475A2B13E4AFFB36665179C5E5C8D752E7356FBC233D290C4AF835AAB0C12B2914EF05E7F947C9CEEC7B1639D62A5547528DFDEE9ECF2106B832D10055B9D11D9E03DA81027C657AB38BCC7B0E96D630E3715AAACC3A530D116805FEC44C4E27F4D09205D11FA6E6DB2B50710EA7627429F44C7C35A24D3DF49B3DB64975F2121F716C6D06CB94ED00DC3A29570E47E0FCFA21CFBED3F2A874778F51C2062C75E4176454436FC5CE68BAFC345298F8B31058079C7F40E248E366CFB4013538F3BFC1F07FE5C0A9A371FDF7DD61C0605F78390B9273841689CDE0A184DCD41B5F3D8A675BE186CD2FF6E7CE4D62CA094CE9230B11C33330503AC00EA65726C480DE7B1827351403D2F598FED8BF3D1CA839368E5EF9030E9808FB28FB4DDE523410BA5D2AD4341EA3F12B447B41BD7F63C9DC429305157F774C7032835123B683AE6DAE1C7A9DCED8B52BFFB1C5A9A66F6F8F0CAE85FB67B602845852F1D6B821237046840E80E2725527BCB2C02540EA8AC6733A0934774D1AE5DEE472D3407187A270FB58DE77AAAE83CD178B9346B21016DD7FDA2D298362BC106068F7E20B610A137FE9ECB6375B7F2C24E7C5361A74D21F7C0E9BF7BB05BB6EF0E960CDCD238F8554EA874B6B300A287139B1D719347BD6D44C855D8E66E29F5F26ECFE843811D79DD1B05E8B392006ECA666035C7BEEA2A33D0ED4799E57FDF45D44D951608F3A33E216230B3F4C6B71D981B80A6E5995DB50C96E64419268F1BB842531972D46DB67C55A990347E13E29895BD213CC7E2CCF7AE8B351B7B48D848A34183DDC55D7AE47A66ADCDF07AB1C9BBA09FFF18C24F275AB891DEDE1111753B8F57EE53E2D364E23AAA57B483E7C4DC95C2FE7FC2B96C6FF8A611157104E52B9E90455FCF307E733AD50AC66879477C7BA84169E25546C699973DDDB3A02D0333E9BFBF165FA858EAEBD41464AC1F9D866BE384F2545CFF20461ECD163174B0E6FC1FBE138ECA496F73C15D8E2BEE8792828A8513DC4919933BDE6E7874D3DFFF89960A204A0CC86CD0222245050675F171CA3149CAB4BD899CFFD044F1C4D038456295DD18D0E13D29B5E25C7B1487CA6ED4BFD86B80ADD50404629A3007BE0BEE425194573C1C77725A07C8B3AC80C9421B2B7994217CD39692D16ED04C31440B8A3D9A13D1C682D412AEB949C5303800D6375272A474FE9D55AA96941E710EE754C10AD44E7D1FA1D67752454BE9A60C07B2EB00CACB09EE2596CF782859083FE26A687646CB0D08B5DCEC8BEB19A429B78C34C6E2C9B87307272BA36D402F12D688721F11733B7DDE19876774CD6A3C4A684F786194A891CB89BE4105D48215D81728472D157852BCED623C80A79CFC3F662E5BC018448BF9863529BC0F80DFBE2F9D347A3D62E9D93B12E45C1219DACDFA61CF628467FC5CBB4F625CE08ED8622942DBF1460A7D764D0CABCB2C9D8DEFD772D19E49BF649C62EAD93AEAAD4F2C5321C1E242AE0A2A06AB71093B2FC7E307AEE3EFF5F8978B795F9FE8D72554CA19354836E4FCEDA74DE36E5AB4C6FAC57C43C79C9F35097DDE6D6C30436146E59132EF2BC690C0F98E651F77DDDF619262953C88D1F692596BC40302034C209D2E05A378D1B31EDC33FF41F4A1AAF128CF1E904A0E1BF685A2D0141A9CE9E5451D344F5068C84BD5C712393249DA2B0B47058773822B66310115D88AD8C3418A2F0E4EBCF9A83806638E7F0BC351C33C5F29D60C1CEBAE39998F7CB3E72560288D1CD670097A083F374E90B61A03275712358AE57FEE017E5BCA11C665C734EF0B88E5092C218FB914D9A398DF2BD890823376D2C26EC81F7DE0491C4F849412795CE7F2BB54ADE9B4B8F20BC0808476589A9EA1E790C675323170F33B148D478C28CA58FE41423C71A8DB160529397C74B61B6E72976211668F547838BF2EDEDCD8DD46873A8F53A65102CBD85A259905B4F124AB775F16387DE165A290DAB10CC6FC614331C8BAB83802399C1E4DA5E9C02521D58F893D84A9B261278EA7F6073A97C0504368A1D87F1EC4FDAD841022E62AEBAAEE30FA25B9E4524448AC6F49AB91133B859DD93A0134023BCE1BE78E4604010827B7B6215A3E39F4E0BEAFA4B389438B7CA9703A5E9C1C8E9D63E92ECCEF656960B5B2C2B233C069C97AF3414DC9E1A62D4C11DFF805CF4125794AAF40E64BDE912F762CF76566D84F86DF471997E1442320061883FCA867B85824D158184B449260D532BFA62F0C4F64251A356A17AB8190B4E37157DF0318AE595527E6AC1205168D7716B757C3604706FB1AC09AA97848E4C2DE2F2AA915EBD576FDC14C202639E449FC5BE5B6925D2447C4FDCF7F7E4BC0D6B55F5EDECD6F7A7A5672153F230A82B9F3A54DF6145E57347BEE03765A7E513BD11A02D69A2B5FDF6F5B5DC7BDA47F9E17D4216075EDAE8EEF5CA483E4E0CCE0364C16D76878F47D6E1FE877B0075C01CC834783CAB045343EF79927A878A74ADD457E4644F8EEB9DAC47E770B33CE859996E79D54801D87ED123C298635D9ED4FC2C1780A995A8C16B2F59738205A50D2623E53C752BA3971919C409691A32E5FAB8FC0C449C10542DEECD979CE6F947CE060896C4346FF7B776AD36B352665D1CA0D9FEEF64953E8B526EB542662041F371B2D4007DB3010788241636FC06531F795EE47EA8881C7E3AA30E3C231266ADAD493DB9CCA1389707ABA584568471BB07EAB9B21520E6B918472499AB99AB0A3B83032B4543E22C9B5DB6A726CC85287EFF9179201E3FC5D70CB18DAEB4DD0174E1EF106A304EBCC0A1F4AC186E8F9D8B60681FA2215CC9F8512C7B65351A105F16F74E7E88B873F6E71F4351F27B42D1FF4958BFB21BD12DB181E2A0F50D7F939C6717C4E4F2C3CDB05664C529F0873F00C6AEB26F9E6333E88A79C1FE02C398CE360419D55C46042114E981499A1FA8E6653E36B401E37F91A9A9A5C3C364C28EA573110182AF2C2FA05FE951C342491DFEC92351C0FA6EBC4C0ACA96B1AF78033F133897D987BEF5B3E46FD908144080E371E2E08E36A0FBE91A6AE4016AA369605D50BEEA02C25AA132D399B8D8DD956DAC9A41131056AC0246E808C95814DE708B5ED4F4AAB05955B0A18EC4676386EF14C59EE805111223F8C282AF175A66E1B0685764346F371EEF17FD748330E3E1E71C8FFA801F2317E599B9538041480FB667B727FE3CEE6C3F537931B6A3355CDDB6B1404266DB2BC3EBDEBC4FB70BAC12AD07037053DF19D68F63E28E78D3083031F9A04058612619B3829CF0776AF59660B2E4079C5A1010D5153CB7AC719B629ADC1DC0A10CDCE1495D7FB6F6807B16D3AA9885432BDD1DB0963F9D27E590F0DB95B3773C20558EA417166007DEB8559D626B75234F551DFB75B0E01AC0736AA54F851CB2FFA99E270BA38B82A12ED31B1A965AC9D61FF104D1B9B6CF8F494595D1BC2C85E95A3EACDCB144707F92AC0A397DDDC68EB8CE09E86FF318C03909012A8653C11D21ACDF3F19926E87BB583FF9C2817100898770DD0419E27F9ECF325A4E6DFF742E21BBA18364239036985F32FD17326277663F4F30E3456B4C2EFE00A9931DFB2CAEA3B0405B81BA0DDD8A5C28B86BFA3653DF9B6CF713B2C66291A53A1F7A0C8CE623C695DDABA40E4FB889744B176939E86FF485D66EE3B93871FE969DDE642470D9183A21EC9D44239458DC569699E54578CD169BE605C5E76727F8731D35D405DF21260D4BECC74D63376E8D8A06E3B7BE2FD6F5368470F83C4B157839CC2783438B0A6793606877D1DBA11E27D73AB35A8A5EE0A8DC08F9B741521420A2A6A1805BB186D3498C9DCF8001415599DB4B2D7FEDC5493F3D8D6F7B3EAD2CF62F34A610FA115C441EA1AAC92A0BA4623396F7738F3A03268480B5A87666C054273BEEBE4D70607615D9DDCEB43D74B3123DD8D2D25DD70AE50A860804E238112315BBE65D94D17860DDDB96F034D1B668C903443297F918CD4A170AFCE3D4CB4A13C7C17352E699B1F4D593D444932F0E98A095A508FE1836E3A8E2F3C6971377D9BB0F3A8041DD5080B28D0DC4DE54E85951FB4D39FADD7DE256921B0DF009FB0CA810D4115B8C33F15ACA09DFB7FCC402E93A456D11C50C097EABF600FDF016D9D59A6038072DE596FC9785A0C855E835CFBE6B7A5904E3650AEACC377992DF9ED809EA2FDC429F341DC98759A726130E0F2482D86DB963E3AE2B2A84A4C0C845B6238573CF6BA87F365C2C26538CE0810A158F0D6D41CB453113973A9E3400831047D393091374162D635486C6E835A4FAD3AEDEBBCD7AAA9D4DA1906EF1E4D5AB0E1D82DB2676AC8EE705309C1AACF4457C5208394E5BF34D8351E932770DBA0DD72B2DA2A3D8469FF1771172122B997C87BCE651DD59B3D1135F1D57CCC733866949C2D43F8E84386DD69448D29D6E6FA2D6096F1662DB840ED1B6853D4A54E7511C7364E895E459319C1858EE4138EE41ABBF5BF4E19C4473410BC44176DC6CD15037D8B384B3A5E5E73A5F0F740C5F2A2E0D9155E33D1337587BBB65C52DBC52C032F82B0FCC13AA5060FC858F34428C116019DEA5F481DE04336828C495ECDAD04581DF323132FCD4D10D483BD4C61B7176B6159FCE5982AA6543FE4A7B4021884EFC9A3C811903C407723B8C7260984B563827B2EEBB0910385B7018047F9BEA8C9FBFAFBDF6A8012048F4F39B9AD508503EB7D6A5EA7C340274487FDBF19E75EA16700310180D43CE3BC3B614D8E09E80AEAB323C3091D1C21385D9382AE259E2389A13BDA51AD32D6AAC5F7DF26ABBB6081B2E7BFD408A1BBA3AB2A61B01AD92370B3D7329DD8D53FE91E1D66515A1D2879EA315D2970D2D52FE3C42F1E19CC1E3CD3202E0C344C5E5063B422152AB3FA234630A5D13663611294AFBC666E93C988DA670E48BF8BCACEDF134CA399D91A5A7C699C70381FC4BF5AFBB9D8A7396F161C24F19CE456B8CB9F6BC04F8EF34F21E4336C55453B56644D4E161521D4E61EA9247431443105DD77D686723425DC48179BAFB0B6B481DCA63AF91D6851068D0A09B0A9AE5E99B3DE3134F2F43B8C04493B3273BC2B6017BAEBCA160A41EDE2D47ED212F2371205FBBCAECF043BEEBBF18860EF7D7CA2EBE81C62A8B8EFE98DFCE21A6B9EECC01245F4B2E74B637E54C80C2388AE527CD1BDFC6D1A6A879DC6F40B833FFDC4C5A5D7B326723E8733749338760BC131AAF46D142FABB027F509988CC03429B1634ED0E087C40637A22D11E2001AF7C1203087173E022EE56CFE57065AE86DF0FC97BB22897E34F2BCC6B25EC7FF1762B2ED774CC7E30F95221A52E5A932297DFFBE10DEA0BEE671674863E0A5087165329D33250A788DD971070E540AE9DAF5411DDC8D260C823DD901C171AA181256988D5B280F9AB714B602E3057466861D885CB0FFFF9E92F22671236BCFAF928009B86DAF50772121B768ABBA9DA3A98217C7612A9F5A61C15227AA3026EF6940231A7376C37E4846FAF72FEF570E408AEC00D4AB5E106D540D6E2AFDC23110E743F5875DB8D10BAF2F15B0F678CA088863A91A8363DFB53123F57C74CD4D593C068B74B2357E1C9BD416E5CB2FD0A50CA693B8062E05ACB0D3E30A476BFF4213F828F15910ABD0714815605BDEB155937111B22F1628380E5A215DF2FEB83933CDEBE01374A7E7B5C2342D982DD2282A9558644E47B366CDD85A67EDA5C08A9ED40327715FE01FCFCC930F505A1E9403568BB6AC484A0AFF9589C856A36751C62EBDC5C96B38AFDBC1A2BCA184FF9EBA426C04DCCF15D05661C0071798CA42795CB8F60CFAAB8042755D741EF5207DCC457D4D78AE8819FE819DFE2ECC9B4A83F55626DDC3598AD623AAB35077D6437EA2136D4CD60EEE838C11260535B3DAAEE12AF5AA104241FA71DCABE96E3854D6E1BE458C6606F0C401B52CD632D69AD53CFF97FF62A382B7B75A47676D5F4ED6F16556025D038E13E572D12853F61516560E547C75DEEA4F4F9319E7C3ECB63D62960E0DE5749DA2EF089FDE59553C3B71F7779DC5D5D3D74F296070B177FD76B4E4A87E4643D8116C8EFD4872E97EE972A62C075642B5D3525AE57789CAB1DA39BE29D64F679D7B773BEEE988FB6314C993A3FD358068E4B242FBEFC3B320CDB4ED6D67F90AAA1E58B43CD53BBD3465FCADBFFC53415AA452F0DD1068BC9D9E93D7215A1C859D75C929047FEB6B036472E337C83861F18ABF2DCC7EA752EF6F15F4D40570072CF78A681D67A4EB2F7A8860F41864AED58F12BC393A848AF6DB7ECD2D5D13061888528A932126E615E3AB7B3C477BA1216D8B24086943207F4D67B4E3913ECF44CC3BA9ED68D023FF6C56642127B6BC03D9A72450E828B435185DFD24952AF690EE8DFAE39980F6BE45A8A268B076E04E669629FE5231CD32F8E4D7D7B2A319CCF8C6A7C67B008B026E9519C27CF9534F9CF907D4A089EC6191E51CCD6F60D6B210B2AD00BE3BFB8DD056FA5D6A9A97C423316D73DBF513821C77C371CC941AF377998A6F5BBF40688B61C0C1624968B1742AFAAEB3758E5881F4EDDEF8A090EA7B7F2035CAC117441DEBDD0703F0BE8E07FFACB0FDF46C18284A5EC55CA547C94A10A91FAA12A17FDFB8E00DE38E0C56E525C0BB49E63F79E3718025E9F4D72048137A2774A4AE4B1F09C1D025A3FCBDA025E7C4901A9B394A3E60321CEDC415CCCBBEEEA4192756A75ED777D361E058F1ED70ADF0425A36AE3A6B3AB914BBFC615AEEFF579DFED05DBA10A806BC679BE45C1953B5D23B1B6E7C45AAC9575A8D46FA9D0DB12FD0C409898425F50DCE60E79F2D39D9DEC916D671440792F9343B4B7461AC0BB8D879977E1925ED821D4EB1058535E853854B1B6E95138901960320963B7D8E1CCD262CE2F4BD9AFF4DFF2DFD0728F5537943989F60D6F23BAEA3C93F1198FD25AAC177ABB5DF2689E530FAC7DB12545CA5C8D8AFB947EE9A82F71A48922D8081D00577D4C285D496BF66D03B81FC27D0847A8F96698BD80EC503774102957161716C4EF9C2265311FD611F5BF9AA3C95E45A68DB0E761E8A77975F94B63FBBA0A84BA14B53BFF093A8AEDACD59A6B90D89ECE433286D639D615520FF21312911DA8FC8BDB327BC1A423E9807722CA2BF94B69BC8F4F7769F11372BB41D7AB1977118932AACB5A5A89C8FD411769597AE8DAE117031FD4E25582B34C2C2B87AF8D7621E6057EECF6227703AFEA3ECC3A5DEEC8297D1D45656928DF8098BC298007248C2713E78C748A068A7BB1044D23926D6E5E21D851BFEAB9E826F491898BAB30458361F46CE8A3EF3B84249CA88EE94E416E07592E23910BC13613D1C742F969DD1ED6B8B2EC67DA58C6BA17CE1C81D10967BB4D724CF0CC0DA570FA93D0AF9DB462C50EEB4318E9FE43ACE3F3241A1E1C0EF5FAE44923F00B7567CE351DA3A75CAC3E847BD435A5322B52007A01CC0B8F3708503805A1146BC581BECE976437C288743D56FEE5DC5AE9C84312B4FE442388ECB722C1AB5519190B8919C15A309BCCC99A1AC4E28227329D53132434ACFA648B8BB3B44A7B3B848E4D3F28C5A8A781E147B229FC661CE77BEC1B9D6C67E6BAC1F81F410F2857408BAEB8A4CFD94FCA1B90336D145EF310F4E2332767872B672B89DC7A83BBA44774DBB27E407B6063EB24503F21F5062F04BC0C10D537F9C19BDE750E17456DE23F940F7F545A9204F36891621CA5A9326CFFA3E04FC9AE104DA44E41317FF30595FFDB4B1EC128FD0DDA073F1EA68A0F0C631B1DBA5379B1D47A77681C62BC1F1B1C321F007B74CFE3A787F9B2FB168ACD24C9F8FB683295AC8F5BAFA37EBCBB83EE773DF48CEA7A64A294A0707EAF007C2573DCBFA6AF84341F0165C5E9D7213590F336E322281464B0B79D98EB80AD06C25085B66FFF58247B5373068ACFF203133FBDCA8D532EA31D1E432B50CDEAA0B731F65F7DAFD24C00C574B45EC4795A97A27526B6EE931E9C4859D68589700A595D2673D23924911B54CB4ADB12B20A0274611A9CF0060799B7D5BDECD92F5BF5BA184ED5F5CB52820396BB725FAAC710DD6A0B04930B6A54D41065C11C9F9255C33C8803DB910595A82C9850830CEFCFC1408D12592483458833D7038331BBA2FFD208F331CCE10250FAD890F16E17975AF409B47BEF7B61045FCEEF346898CD260760B80BB9AA7CF2760CE44101F7E077FA75445CEA7429E6DB85917FEA8839FD2912605BAAC1F05487AE7AB4A76BAA8E9913CC226B7B9224660AD6F88F1E08A4DE9E99FE10FD3F52988978D1B4E8936B7D2F406A5F974FB418072035214F7088CFCF693608E2976ACD079411E7E90AD7436FBA1987C4E56BB30A97297BABD8D96B41164F2FD4AF5A43398E7D32E8401F15B5997EF6F13CA21D0EDFD5BFBA1B2787D52661BF0A5AFABAC16FF3B27FDF4E23'
			},
		]
	},
	SiggenGroupItem{
		tgid:               10
		testtype:           'AFT'
		parameterset:       'SLH-DSA-SHAKE-192f'
		deterministic:      true
		signatureinterface: 'external'
		prehash:            'prehash'
		tests:              [
			SiggenCaseItem{
				tcid:      84
				deferred:  false
				sk:        'A84AD3150675B6DF30E471C01D4A88230DE36B71544E4B5778981D4473A5804C93F54398362F1D164D55CAFC162545889C98AD42A206FD335911CC452CCCA601838EED5505DC7B3905F028F173EDDD0E9C99C2A01C1B341C65114F3B1BF41408'
				pk:        '9C98AD42A206FD335911CC452CCCA601838EED5505DC7B3905F028F173EDDD0E9C99C2A01C1B341C65114F3B1BF41408'
				message:   '7A17F43ECA4F29A788C35E8459490E2F79188043FE0A339E7952B5E11DD59D8E8CB51199837853EE456E23F87F3331B94BBEAA23CD88518CB177B61E3E6F15ACBCDEB78B025AED243B4DCB5096E4162F70F4503381596C444014F3719C8E3C10BEBADC9663A2AD9BF12C7C3ACC91A0A4E853AC7B7FD46698751A2DAFF6DF50B88898E13789FF821D6FD008E7F1E25F6EC4E950ED47C5A9A0F16596E6C01D6CFA146E1D2C00658E3940F441297557FD0B01EDCC62D96426A5C4E29C1739C311B0F97D3FEFED605C914B2A516D6B6E828D7CCFA9D2CD6577535D0A8C5CF6DA649261AC97F7E57ADBAABF9AC751B884B0513E93F19E55735D9075246AC80B1C2C137C0AF21BBFC1206E6DFE452AF6EC78C8D3977822EDE09C53C856B905E948A905C5BD3E304C84E9B7B6DF7FF1C725E72E2A5311B421F1D0BA3A3E9FA879D64DECEF0C50DD1BA31BE44C9A14BE9BD69267FF32DC36359912159B5AD368683552CA9D1AC75A8DE761078A464D34076B150EA708DECBA1EB07B766DDC47DAAA52B99CE1C2AB1E43970DDFE7E223C5179F35FD87D0E94CF20E7C7CCAC93FEC56085AC839EADFACBED8CB59DADEC88B3D364FADB89DE2F52AE387C17F69F70EF0E8BEA07D510B574CEE9B6AD6043079CFEBD6B1D830C504A8C81945421C9B5A43916E0B48987713F827EE7DA28BBD4438C9DE0AB43AA05EF40738E465038F2B6C4DF693586933ADF69AEC889FB90BE1AC8E48C137F7A83A24B6748C366DAEE4A07E26BE6D69C2718B15F26C64D51568837F5213E82F9992FC640D1ADACEB3E8F7515DA5119F50FE9220F0D18A949E31D15F5AFA56A6360E13485DCE6864927BE78D00F306E6B7EE69A8BA1E2DBCDB4A22657F7D4AAB75F854549BD98DBAA75C3F1E8E65EEB0A750CCA5A5CCAE8A62BF11DB791FB0D19A75E2EFB3AE4784840F6568A8806BFD25AB85305EE52158E81802D35E11CA1CB4E7AEFA53045C2C811B8AC725969265826FED332C75B9496045F41FCAD8901EC69B0F3AF5FE6D02EEA1A6083E81AEEC27DDABFE2080A7C422A4E8C0174ACE3723B958C482CA333E6E1DC3C439DBEE59061B5A990FC3D81F5F8205292CCB20A275DFE41CDAA5078266BBB208AFF74627CE158B37ED441717D623798A4CA9EA201673CB7003BC6E915347ED16EBBE42C90C41D316EB4726415FE7D949465ACA43C2ADB6F2C05279913C767F1385670FAF7CBFD516FDBCCDDD668BC27D5D9B17C25B628DFB5DCF88D168C0D3A9149CDD226526D45E2D25B6509914B24933D262002F93A0529964D6511DF24CA40D56E228D4F65FBF9B37660BC51750341096D3B564E10006B5A228B4E67F9583318B77F948C2E00787C6E13FAA5604C229BCC0B3857E2F75403AEBB50DD7868C670051C9E979E0E14A5923945650419167369C6CFC0C938345517329A43A50BB6B478FEBF76BF8B629CCB0190174D6B3649FFF6E92E1C3F6FC4935D2300AAE0A7235093D13A63156952F5EC0038FDC8B23A3345234D2E07474A38228C28DE5789CB3A8DDF00A6698E234318356489A8E72085015734ACE1B1309377A4F239AC6B2B5089E0E4E8383B8B79D02EDF37DAC1DC14C6D44982DA551B72C838E2F508F372F86D3F4B84FBE65A4BDA0E01FD23F9CC5A99FA2C1E639890D565E0CF93876588D12C0331A61B760FF3F3AD1B6A2A815397CC695A91C59EFC9FE667FB0BD94EF8F5782C7E779198C3F48BF2BC6038763C60EBA8E27F5B01FEAA7BC23FDF6A9BE5B00D53E067E23F40AEE9B692C4497761254665A6BFFE0649599461B6D146ACAA1EB606D79A9B83C69267E086A55A920C3194868C15B99CB6E5ED7BEBA8D1A88F705BEC5655A9F6ABD37A5F5BB5EC37D57F0A877AD61D060B0D5B8090465641F1C29573DC2F1216B90E5CA91CC4A911667EC242EAC36B25E3381C696B6205077C972304C652B598C1F44AE5FB003F2776C6E3954ED3D815C75CC692C8D30A04F457A95BEC20D849141115C2D83381A9CBE43C7666F95F26F210259F9CCAA9D7B723187DA90A0CB33D498FADF9CA25EDFC625D71ABC1270DD45366F9D41593A4BF0F8DFE207D0C2856E8388E0733795809F9B4306E68E6442139FBB532639B75D896E173232EE6B193CBDA92064946CF08985C708A6C3AA182B02D072E9FF3307A3ED74D0382F166693F9CA90969F54E412A54269416B3B0E4E5F5149450F02F75E4FBFC9887FA5DBFF1863E1C1F8677C5C2581FCF6915753A70D5FDE0B057F07EB9C990E1BB1199492490A98CEE20BAE3D5C5EC416FE93E75DCB7A92144824F9A122D3DDA6A4D8BAE998EB8A78A52F219F7416200F102ABF6A3FB2E46BF32D8DC3733DEE03AB12537C6DD431AE0E1700AFE68541C5E87CEF10D788B9084518BDDA99889FB5DF0824B5EC088BFF3B96F2F8BB2984B108275C12F3BD1BDFD84F84E9D37D44F11FCBD96B3649FD349FD2CDF3588147C9F29157EE89AF71A8636AFFE94D1BD2098A4B8A02F387425015D5C265558F3AD838C1F5A586DF3C99DECCE2889A031A524823728369809BF846DEBDB649407555E399FC576E1A2D0CDEE3838F7F892EC39C0BB5DAD51E62252963CFA3DC1B7D625C5201C8D6A66DFDFE57A1CBA5B55C067299D1B6A2C1B7F552C30DDC182B5470AF3944CB8FA15D6DC2689C9D03C4F8273FD7CF308C2C9B912D916A340420668AE4B590ADDC8BEE41CA6DE34E52D586CD07020C7EA639364FE711577DF327CBA5B6EF629A820F393C567579C26C82B2750F5D5BCFD61D7A575022AD15C834C734204FC1055A962A62D1D29C2090866284371FB2BA6BEBF577F4CD30BC620B1EF2A60A48CF06E994C217B7BBDB957F1480DF0F10E7376D3E791ED7EEFF58321A9DBE319FA50731934806EA27AA55045FE3BC88FE7C98CD2435AF5000AA319BAC3F5210DFF552C109CD8BB9B45BA2EDC91F82108B04717CAE8E26E27610FF2F01BB35CA882E23D204478D6FF9475B4B282570FFC93356E209EA3F03D75708973D84F10FA6CB033A1F5B53E1E68B66ED91FE498EB82CA402CAEC959B68332D582973FB5024ED4971A4292C7D4611CEAF85A73704BF321B28D525FCE04CA7634BC899F3A52AEC84C8F308B0C3558928B7DCD242DB7EE5F21D29264CA9B64C7A54FC81F66EC99B81D872B5EAB15F344F21DFB33CC70C5FCDBF08CD40BCB4F78EEDBA0FF7A4AB086B09A94F2B3CA50AEA69D301A1352A3454F426A17734A52B17ADF29FBC39AE123370E8670B6143E4507001E5D7DC95717D763995C6DE895360A4B07F20F57AEC5FAAEE46A6A7BA9E89ED8FF09805CFD81D13953715FDCD11C79F0EB5FFDDD1D06099FB97A4B28502BD5F9383F040F27F6AA05CF2D5EB765B4292F93BBA67EE2D7170318A852A787A166B228C590FA4C0DAC92DEE0B4340A21470C22D3CAB7DDFEBEC939501CD38888E6836268D9ADC14B035E73837CA1A05054347BDB306D24C91A027252464F6B1F165A8254855E56C3E75340EF80F800311B7F9F88F39EE368D8E8C72F70A89F434DF37B7CD2BCD0F4BD6F7914D5FDB1E232E3FBE592B81392D7541056521332616716EC32DA3214166532400630BABCE93E1A43A30A0659392556AFE6D33527FD75AACE92E6EFFC758605ECECF239E8863BE48B7911A80C36A8D221D6A89A1C511F323F1941F8CDC993554C163D020B472D5781EF864630B5C4108AB3B990CAD21C29EFFD8116DEBDD312C0425ED0473385DB67736D397B0E30C12F1FB5A1DB5497AAE78436912394CAEF2802556176F42F405495E4627C04AE258FA4AAA8ACFC1415A3D4C47774DA714BD5EA3D2933C065DAC7629EF06A3B7FACFBAA6C94E09FD9662C8921DCCEF7A3F2854E9DFBB0AACFFB388B488662409EC5B1936E17CDF69A73E6EDD403BC9E6510E800300800303F6AC1398B7B13BF53008CDE7A34088BF3B6579E2CEF149135C4065B45B6402BA32BC777A3C0ADF21112DDE894F2626C6B2EB77133A45C06E165FA386D25D130E921D0DDA073B9AB288B4388F6F6F630FC738017E7294C740967EB5D6CD57D559AD3DF8B225FDFEC459E9B7F18656ECCC2660EEA7A6B04C8ACF23C8060FF49C30B5CED64C2B8970B5EFA83EBF2F86645E74B5CB59988B18737A244B96B3EE7C8898D787FAA55171E1CA8732BF33C6AF0ACA8BE47C7D35183DB98BADAD7B3B4D12676275CE912EDA6922389EB0B8D1FF27C1B6D1F100D3FB1EA619298FCAA42A5937EB9132EE60C19C7CE5507843BE56E31B68419594750E08A5543F52CB575E72B0E26F1FB50A80135C66760EEC9072D57BE4E71926DB4BA70B464D7E842E02F2F43D08B693C2C7F2717870D02C094EE2C2C380CE4A52BFB9A902D28D0D018BCD46A2182B734598FCB3216BD694E4B9EDC34A701FFB59951C688C0C3CCF8B23ED4F05B4D5E7122D42D37C27DF6F1845A53FA20820FEDAD30B880F4DA0887C68DB00DAEEDA89F98FDB6B7EEACE551D1BA63C84A9386624B82DD04EDF76ED98B1BE3A7CEC8ABE7229E8DA6E55B6F8B34A57763B494A3AA357FD559D4CB3D26A49B125E371AF6491D175DED3DBBE221DCB2CF2A1D13759E791BC1C511C8FE808CCB62C77C4C3D03D094762A321DC5F644E622D34BCAF107638EAA741DC6DE9341900A02B22608FF851BF50E1AD82C2390DF8BEF5C401097CD15ED844BC21FC5A390025F4055D6D0D67F135C62BE1C5012F5373D8C812444EF4B5888F6DE7E997758CD36293F19C71C1770818400E3269DE462C95B961D70C62C9E5A1DF2E74700985C46E5B93575BF93D3A9F1EB708EA6757BDE257E31D49EB2F05EB5D85BF0C1626CF58E8A9B19C288488D6ABC22B78B533278E2A9A96C8DEBD081D3F8FE07203E6514A2FCE2D9EE5E87CFEBBFBF6E33C356B3E07C2E27760EF170638A774A57334C292A567AE20612F411D0207B7F5B330B4B42553B6D68906B1CDEE8EBE36F57EF663E1AA13E0E99081BE996B7E12BCF594F6DE7A2469A8B44CC95897B0F2EDEA88701A74FB5827832E49CD6F8AD5C00A659F81AC117DFF10D8DD024B7417EA4F1E24313E2D12952692FFF8138A81915F04CCAF9B420C0EB9BE4787807EBA73265D47E11C24D4D7053AC3A82037AD58606D7105F73E37970F306602F417DFFA3B103FB0D2F1FED00AC3DDD2D90B4F2FC13BAF6068F593561E1AD31AF4DF9AD31DACB37F677E941FDDE9FB8A8455A1E25B6AE28EFAED96FE8F973F6701CCBA064E62388AED9A8AB3CAAA5E0FF422FD5D81D4E7BEE5E9454637A119E2225EBA2BE9FFAD71A333C73319C8783033CE9F997951C5BBF8A3F5FBE3EBBEB4DD947C32DA81DE83CC66AF4790D052DBD52931F655E786AE9194BDB87379E8527B58136CA45D5965C4F5810FF05750A66C7965CC3E3A0CF101208033F793794D66AF9EE186BF554AF5602062E887CF11D8B54BFCC75EF20A499A2C09985ED5E5587987CF79295BB8762D2B3034569B3D3A2882DD78D1C6FE7F081AD267CB78109054B973B4F94A6B82C4CE8E5D6112547C93D5107F764A11FD4CC8B384DE7D34BB88A156BB07C10F48F243B2E3B44B37CB9FB0E50023A931BB748B8608835DC677B23298A8DDF42D78D54418A7F58678C2C146E294F4F6EE114A24BF3539E48D1AEBA87A3D0E09027255D9F711CA8BD023B0CFED0068B2202C6FA6B1E0767352DC65D333D5BA3982BE575B5715135DC80C1525A89CB0E2EE2F7E247690B769DDACFF1A7F8297F559695CADF356D1AE40D637794A442041F6D555CBCB03A2DF5C4AA228C35433FF856F79D8DEA7C833EB4928197013A47FD5B27EB3721D64C3422B55BB8ACCE778FFA78CFEC3F6046588D7D93FD6E50AA2063CF5AADD33A7026E4DCED31D410BC4790F0E7AB5AABCCB6D4BE7291FC311010E630C968160880E2232A970C161A17FF0F8F2E7F6090502D3771B5531C94507BE8044CEC0FCBD7BF6F483BAAD804278A128E254CACF914321CD933EDC7F02A5FD56F103DA5298D35DCDB7875C36C066B5E7D4347F325EBF941F1159D00B39BE8BDFE17DE6F850756D6197298F25624317734A162D8E85EEC4E80C3AC7F644E4F746BCBE79E7D9FFFDF1C3051123A79059E95024F020F5389E5B55C0F85E773076B84D36B5BC2C77983A4722C7244A1AB8F4994F36BBAD347D626A965F723A45249A296B3E6084E32886D09D6572AAF8F1B53332A39BCA90138B974A9F550E78D7BC95621D3BCFFC273CEAF15BC0C004BD09FB6DEB11F1CA0C46970E5CBC2013883C5E35875802FD132E449565C6E6BA99E406CF7896A535E22CCA2038E31A7BC240C8327B59F8B3C963F48047D3E6C666DFE17737F264507ED98F800BCC5107BE8C694C9D5D8A7B5B3EB1DCE7141F61ACC5FC89EAC8F83B9D559005D553F27B30DBA45745839C6359DC40302DF1A60EEF54D40E4791E352E3AED029B0E457AB6EEFCE9D12FEC680D4342BDE2BEBEA7D7F50EA2CFF616B0F78C7460C04609785AA6C1C186F255FC981D36FA2A15C1A29BAE48A5869F2078AF83DC272C8585433E6CD2A3605A55209A9542F06EC534D3B3A0E6468948E42D4A221BDC13F092DB0EA4C05EE9754381F4D2EE6BCD6B9ACA5FEF17BE6093E7FFCBBB19A4DB4AF288000F5B089094C3CB5F46DA7147AFE963C6F726067893EB69AD50F2AC40A2C8CE43351BB6CE61C186F590524BFD944FBD685947A31936BE1CC62A69521AB85BB192D7'
				context:   '53AF0E907296E3BC83453CCA80085C3B02E551F004A1FC57FB622BE200ED01A29BA906879DDF78863A193D06155E7744CCA6C6C8DCD9225A37AB6FEB1D1ED5C04B5228F84D28E2C8AD2DCA26FC33026B4D4800D5AE4CF4C3A154B07FA725B4043F393918C9C58DCD7B7414D09DC3AEE72B1710D12214FA856AF2BDDAF55D3DC1FE67EAAB1B2E825E1A23EAA8D15FB55E2FA6DDE5E7B26C2AE455464B23A7F0661CE62F5322DE8E08FCF8848F3FDFDAB13DE182E6C35AA82EBB0D89A9377E569EB32987AC10F340B18DA13F8FE127376EFE7DCA7A45A48FA492404762901BAA3B8865B7764DD92F085BC88A53FE3A6E026F19C4E1B9DE036AA0D5853FFB9B'
				hashalg:   'SHA3-224'
				signature: '423009D1B28F66B396101A443CAEB946BB96CD3A3D04DD07BCD2663B244C20C381957BEC9A27E5F7E521D67CA1B22E9400F535414AF196D6BFDB453032C52635035A45E2F128889460047CD8FFAEDD42E3214F48330F7E43A56C885B97D82279ACF489E40526F1277C42EF96FC3FB99C961490319D3617D4B624D7AC6E55A94791491273160F967DEC2C859D12601F0A6CC2E970EC23F7DB2952C7E28F183D96C911BAE220D336EFDD1F7C1E6CB48F5BC9BAA029D95A7CFD9C9BCF325C7766B30F473057450AAC22DC68067299E46C025D4A2DFACD0F39E26036766B3BC4BEFA536F97723EBEF3757033521739F1FAA532C988CF9AC618BCA24489DD98527342EAC3066E7C2B0750A1D10C285CE8BFF6E98AE50C3C9D88A1E4938AB46928BFCED26B46BA2F6F6D84D768C846C02AC60523A5282C29658DEF7E98E78AB6F9CDE4AB86C2B9204EAA670569931BA878D71D4D61B78A150E7D4AF3E51913693114E0E77539B22C433CB2B74CCE68312361459426A003F33AC7846200849CA8AB326516E2797517F0A0242919C24B20B6B34D126BE43A5EB7206DFE9AE06249ADE1E751A4B25A6E32E98D18DF7FDE2C5D965D261BC747423CD94C86C4E707DA01CE48B7F811E28BD3519BA0C5438DE51AD77FACC56F9F31ED899CFDFFB18463D02C0B91DED66FA4003E660089AD25E006F5AB19CC05368200536D70F161B45172B5D697D34C0B1C465C90CAD04768FB8B22A337102E6C8DDE68FC82155E97BBF95851A3320DFB8DE4BD9A43EE333C7DFE701A4ED42D8CAE289EE5901F6DC33679A62602464293AEE1D357294298DAB3126C40AA1681C24A4713FEF90F76A9D98D71C8149CFD9226F4EA1937BD348E1DA43D17F31AA9BBC647C5C236030FFD7EE10BC6C80F3A810A9AE156C19E1035BBD0EBD9BC8149726C7C416C86532FA33F00DAB446652E02F556A1BC27EEAB8F3638DF6807C5CFB3505518B098E2A3B6FF3817752E8CE02A50D84F253F73D913B1A866208AA2F258EDB3AB66269BD3DEE7E9254CF44F9FCEF3D8DF427726E727913503349C2C574E3129A1F4485D5A550A6B0BB648B47AEA75EC721E5509C9CC54B8DF9A2070EEC9953E431140BD216007ED695B9607B3CEBE947B1B7E2865F523AE94D3FC53894975C806F1E271EB33AE55D24AA4E1FEE32ECFC2BAB1069B82109F6D89FACAB730375F2438655F8A592133F11FE1A222C484241E75BEAC11A1676382B7F4ABD7A60DEDDC1E5F55E913E4F136A3785C866B0DC0444BE2203AF0CEAC671B6FDC6A11ADED63E9AF766518E76AF99BB417B4884C2B3E63CF3EC7FC0C50071413994BE0731432FA78239876772206EBFA9981152DE59CEA8C960380D453B55733ABD243661E3E89FD972EC7EF1A913FF4687D132B615C8C85B8D4742B012F0D775ED2D46251B80C1A669101900750492AFA53C48FBB47AC0812AC52E4978298C9BF363CB83432EFCB8372A6FD47FB216D499B6C9E69248461FF688CD1D6DDFC6CED83D57ABD51A56A1DDB663604B705E5D3B02148AD4984E4DDDBB822532CE5BD74A3ECFF461508B03398ED8CD95FE9A5CD40BCB61DB69B85710C885E8A93AD8816FEC8C9EB553DA003506B3064A3484BA356C05E896469133557A58122DF84D7C8E68E7D3F94B917A5C9EA305A39FBCFB24A6C4E3026383A1CA8BFF92FFA50725D27E1AF029B45A3A8495C95F5A0EE5371D48BBC4A7EBDDEB6634D554E369EB7008592364CF64F826A99E015BED20EE08782D35D12203FBEBCB2DB181F66CC7CC7B62EB8740764DE4C802157130EB51570BFA814AB6E70674692913A00FE5FBF0A7F341E1760D2E17211DA3792F3F7F0CE288CABC3EF354F4E807E7A0A4636BBBCF078B558C770BE5AB339ED018BD4D96207DFE9C37B16345A8E022AEA4C8E903315ACB37B1D95DE9CF360DAF641005F794777A73B2217372612612EC660CC09CF8E0EEFE2487B37E374808AE07488154DB1C83DDF3D7292A98305769875499D322E4A7C766DEF301E6FD5927511A7EEB419ED7FD6D978D795246F955F8B1077C71C5564605F423EC8BB6D4A359AC5DD6053F97DBE86F9856FD20308C3147075BB9D65C7D858E87224897360E8F3F0B16CCA6942DE477C74761834CCCB07CC2E9895E5B4F7FCA085A9235486B195D5C29B6295A945D3EF9AD1256968F845C4273270E1B068496858809486326A0C4AD11A256339529765F2FFEA45B976DB34C4147F27616790A97A7E13160E6938E1246ED502C15968D6FB64434C7B0A567BAC387C17CBBBCC36891F8002806DE0C96E78041EA89710BC237533278EE8221C64104CD744B30B5121254D5BFD559135FE718A5CCB7A35A211EB3FB9CFA69348A52148FB65BD89A438BF161CA21B82341466E34C77D14F73741A007EF649FF2D0E1405CD25C947FF87F27574308AA66396655087D0DDAEBC8FE056C230F1A37EBFF4A6FB05D2D9E7534380D1F74817FA05A0AC616D5157EF605F62DE6101F969881DFFF40AD81EEDBD9FA2D455FC0498E203102C875130B9D19CAEDBE39BA0D34503BA02CCE916C260AD69A068764B36AFDE0B6FEDD66BD20C249856016FA973E5FDEDEE3AC49B985D4174AE25BD5943EA637AFD8E08A9823A75D8761B50AD9AB49E9A3050DE0F4E59D07B675B079D6A05815942B4713832575B7C39B3B8BED85EBDABB7CE08D183607A8575207F1E07F6FF245B9C6554DA8F8B618934DC9F9C4290D0344C11227E07906726B2527837C0C9DB75A530D9D361B3B2966FAB43CA7E1F4908466A74E62CBBE23DE564EB69F3D635B5CC291BE5CBBEB6D3161F7DECB1A79AEC55C83E37097BDB7BA35ACA22B92628B770B6076BBFB992026532BF0E42C3CFCD610EFF88056BDD9D03722BF38557B221445249F504A7371F5CA880E3B7750383258C8E1B4D4943B68F601F9E216EC6F80E3AE77E9817D35F2B150CB5F8BB3B0FB3F9F89689C18C8DE30FB30621EE25CD2352BB6934DE765B79086FD8B69C6DC065EFBE11549D95D034DBE99FB3379383647289E45CC14C06E340D286BBF8D41EC15CFBDF95BE720E3157F2D8FB6740FF86109F73AF4CF4C05EF42035870A534D50CCB79FA66D0AB0C0F51D5FC86018C4195DAC748910DCD51844AB41E88592841DC452BBD6C205A47E6FB0D5A85D688AA744C770A146D3734B4DE95AFBFBC03E6972CEAD2AAA3F5349E2766E7798BE122E1540769446F25D59114FE71EFB9F7602A3C589761B69B011FDE928694DCB2219B06A0C2A8D72F14F3055556E1DBEC0C35227B43F03398993DCD8662D0EC80ABE4CCE1ED8B390301B463DD482BFAD17699957100BA4781AF4A8B258614064C8A755884E6CE2084FE1B8D03A82DE355700D67B77E22F588405018A489D7775E03A8E3460FBE86A23CBF97B3BE94E6C166C865F92869DB6AF226D4BB7D3B5014A3ECB6C5CA4D8261830AAFD8A18ADE01E360B75F12C57B7517559AEF14E2A263442223E4CA5C759C21CB13A6FE390BDB39B922DAA47C36F70863EFC0A9532252D081B5F1FB5E6FD1738561777053F93EE569EA47EC3C7166F9630D1F310083640A9307AC9BF8E64F93B11AEE392E46A0BBFF30DE17AAAB16016A8660DB6F0071A7A894E4512BC0BDD5831A491CF966B38F718775BBA9900137E2A3B5FCA4A2758FE60526838AA1D2109CD8B34702B2284B63F2594C0FCE155F44B1E40013C3C1B67E308A3B68A2E5D7CDE30390A884D5E15FEFBF21B5B196C14592800496F0E54668B4F474C3FA0E6C04DEFE169F590499DF5F8CF6930B7EA7556BCDDC5C99D2CF165D6FB90DE42A27985383EA310C64A89B77B08AF8BA552D82D68EDA8238B98075968D322A15518B1A00948A9A029A8FBA3DEC2710698A07100FEFD3BF4FB2CF1A7899BC58A8B3F6AC75B2EB0C1E23FAC63638AFC43FFA2420B920BF6430C84567B9150D70774CCF264F197BF2FCE70E65E7E9C72D899B8772EDCD709FFC5CFB2D24F870CF8AD8984485B80122BF148E58DDC3392C8A02B90107754E9049E085C969B4D53D13480A0EA8A0E209C5FAF9BD3120AE502EC5A9FA22AE0F6DC7E7D2980539CD2FD30BC19EEA79836109220F734A68EA478DEE1A30FE3AC69723D7695A557479B56A84743AA3065182982A017E76CD197611CBA67EEF8E36744A9A64F524AAAFA800DA58D64003606DFC21D0A5E42D5D9A96870D69431F356D4F385FFA07374F33A4342A84A3E6F12D7E1CF52941A78F37C02C938BEA17638335F53829DF811CBF3D86C194E1E3807F29A4A6C81D7A38CBEB533B3347C07D610F95ED5546C598F5169FB80D83B9EAF1D0F4C631FA1A4E84ABA7BA0B29FD12F3B8C838493097E2A8A430C48EF6D66837B838E22295E22D8344BC0F1DD7CCB7B9ECB67BA12056D979271CB72D87A682D102AED25179E7774586453F5BFD968816E6FB7DC8A343904B82E4EAE052E4A4F1A5C983E4FF8B9EAC658DD3EBD647EDA6F73ACB9CCEC72D1768553F3430C511C3AFE48435D06310FF5B1389F5D8899A0565BF44A7D28E9FAF0B893D8412D3B37B132A6E8DDB5F8CC5A0D97DE271B7D3AA194604C0AAE6056730F1D26654BAEDFC23142384C8C2D12A3F36AA2C03DE01B1425CA32C0A1B6D02A0B7F4F02C27DE6FFAC02E3A7A22AFF050D2D0E5F0936EFF122CA0D7A1B428B0267DE66635FEAD2F4D2B54D0FDF6CB2C1289712FF041E49031DCCA0F006E608BDC332FB2D89077FEC4BB644B904092C53C42007B5FFDD92A210EF2F14C41BEA8FC22DA94D7B516ED0A1E199DA43F6C01D955D662EF5F963DA19F7CDDBF8FE88417A5E8C0B50747F3932E3D770E8AF7706CEACCE00B1A8B6DEC284DCBDE34B4D44C557C9E912FEF04EF9A87DB53FF1EB961A15B1D0F378E9D2A405391627D7CAA9B2A7F3141DCEBC18A84757E466F82BD6F3DE7308A76A2FE923E6D8C920E1E4DC1C45C745610F3B3ADBEE29E0A1695AA98E1B66F787AD662D9681480EE45926A783ADF122F1707750773A46E989CBDC1E31CD3AF8D41F30A8D3DA4642AFD895542DDE184C27D206C41ACEBC482AF30F1414AC0C9CC57ACDD72A81DA63D391BE0945C8C82521067632EFBF0C964F3774A31A71FD449CE199235F3096BFD93BDB06F40037875B253FA42710048B37C04DF25D24A25B78B05071424471304A3BE574919384FEA342B3E0D8AF062523A48A542306A1DD9A5E501285A92744911C5D6118D15DE9AFCB64187112EC15843999F56DEA95CE10D4E79DA9A1C198E003757FAFD04B6472D2D2A1FAE5B33CB6D7D5954D5A4450E362B509D9417CA478CA0F1C5932AA3CB5C59B01EC6B8AF132B8783AA62BB57E1D3A720770CE060807B9FEEB152C7E918C4DA9FD9B0DA98D3CF6C45BD6A484104DA179236CDD3D4650E027F9A82A3DF69EF32526D98D9A54A0F27CF02EC78CE697DBDFEFB7634A8212ED010746EEF1B72A7A16BBEBE82BC89E14D00C3BC01F5E1E859B3029DA4FCBA060235063D1130D5FBA5398CBAA14BDCC0978AE3B27DA360E020A313BA1166C1E38C3A4C70703E7EF049D6626EFEE054ED43BD983033E0B4D3F9383CF649E22D23D870A71AD3310E94F8C7CC34F9691BFFCD547C1063C506EED3FDD4516D555DB2140DC281700D36EB8B2EA9F45EB6466EB4E42C7870EE475FFC4520A5511471FACC257DD52EA75EC9EA6C9F0741063C29F7457156A3D602C343A02F4A2DECF7E141C0BFD1AFD9EEB0C2DFFDDE94AE448D7B34D9EB0DB331AF01F68641AE25707F2AAA2996D931CDCCA4DA2F8E21739A1B0AE1C7B11E38B47F4E20036A6FBEE22B90DAA4669AA97CACAEB6137CF9C53F1AC965F51D0C51E97E87A15FCB6DA1F752C0429D297576CC096487AE420C936428E2D4A83883D2C57E7736713550F82461617210DBFA214D7C948F0FEE87968F53F1896D979DCB9153765ACA71CFD7062B92584EA090D9C195B0F476D849385A642AEC6F2E7D76698673D611AFF0404DD2495230747AB90601B9A1200BB3427E311E0086EFADB11803A8B365132A6200F1105D2FECA7135E9852D5805EEA2BA52745E87B897BB4B4BA5F0790A39FB33E27573FC742B43931FABEB34647151614ACDEFCEE224909F72FC197ACBC3C13FCE0E5061AE53BDBD8BA9329BA6F3E0BF58942B38E3D5273BE105F3EEEB4464A60548396624B680B3C576750C7F7C9D118F785C35B9DB010B85528939B1B32E1B00E35BC0B92785D390C2098B50A188EFE891AD304736EA130D88E0B7CDF55073C6103ED5F5D148A9F4FD0FA89AD10916EF61BEC658E4CB1C7766D1056C817F04546FDA5B075D8B43B9911A3055EEE1791F9DDD4422F2478A869F80B13B8DA7169FC2AC4B6AC72E190F3E93ED95D411D4F2485A0A02B1DBD7D9DF98A305375A224163D1B56322A359D58A0EF7C2D34A8C3901455F20E216E55078DDBD8F5D2F1882D4256B6B4218153903B29B82EA20E74DD57A629AAA26557582E1FDA861AD65AFF571D032A7DE43768C8DC28ECD2ECFAD8B54DC4F3B5D8D6B56B3795531A94E7D7AE39CBE6FC5515B6FDBDCDA70FF73C22A158FDD487A13E8445BF446ED3098ECF2FC825ED414AF417EA4E3B1EAA5DF8DD37DE49246964C62AB354E17D16BA1B4D3B9FD22F80F19462354C2F408A127AA28DB5A5A67FE0069B5BF1E6658FEE91D8F28EE815D88F20F224F0017E8A969B130F1CF57FFF296451DCDED65C50AB87C1BE337E2705339E91637A6D73E49E1E7D57D0F38A92A7167101383180792846AAD13B49A57048E260EF849B25E918844A4307E132D976B1F5C480F6E927BEC73DFC588460CF02A7906CB527F186FF8B2DD3DCBB0224E7242E2B24853E1B0F9DE528F9E3A325DA77FDFE04E86A93C504B04A74A1FFD2CFFB98D2D38DD08EEBF8C2F03958138E874313986B311D63E2EC399B48756711B95BB7A4C7A60C24DDCC4E59A302F9E507CF46838E405D8B36B5AF45C2837691888BD425558B65EF54D0EDD203D473FB6729FCE0D8283F8F397E4D6F27F87057029A401503B8DF0F722AB30889839B40FF69191B491BD9CAADABF0F9B226A09957D6805AB0AFFD81568EF9E021BD7B3A9167B48D1224B144A1D6F1BAA8A8EBAC5CD6F9F38DF97694948FF482117D0FE5E6996442CCCB392ADACE3707ED1800E461C57EA7A3783D6A01D6D0FF31BCB485C18688A31F40AC08689CD182FA59377B80363037CFACC47BF2A4E38635348485D8AF1D41D40FF16FF8C4D5DEAC62BB45B78FA3DBA57F1C9F9A25AD167DD9EEA855BC2E432791B4C36EC538C76C3493FD6B68CE1B9829C2A653669EC9D6063B9D9234B43B70FF6DD5AC882CB5A74912C3B3C8A1D86CC6316C30BA97F6D23BC171B507D18C8EF9D799FF40CCFE682FAC499F3C1A94C2C4399E6B8915DDE166E71E1096AB002C60F8EE398253EBB0D7F5E111E7F606EF8ADF60C8BB56E96F72639E5BC2AA0D3A46748B3D8FA361E673F032B540CABA3F09738D373F64DFF3BB382998B07B0F535C1D05BE6FC7A60D818D06A10725F993C29C1FCAF8D6ADE036F0C33D3E07925024AE49FE0E4B3E310FBB18D825E59E816A5A842CC46CCA4B507B84711F31C42625983C6F2DBDEB04BD905736792B20CC5AE3EFEC4D1D465FD5F79C785AF4B142D31E6269BA4170A2D59F5F0170E875CA2547362BDC2A0758EADD83A1778DAAFFA07ECE222D7528EE815515F5C7982CDDC08C9804B6B49CA75E37000E3E1603E4EDE66B208D4061FDCA5C4FD944F1D84BC0F2885B6D819973827A37AD6BFC9FC17881CB85C1C216608729F8C3AB1019224C96DB760A7A54063381B18B30178C4193611A6632C3A00E89D3ED1298280D28D5562629B9CFDA31FB5CA1D3205EAF89F377C6D44F60BEE9D066925D7C90A657E6F3B9679EA5D09929970B2B975FD33A4ED1FA83325859EAEF6B95E48157D9158F0673A9823589766E31CF08FCB644B173BCCC5E469748BE71625343B9B00BD70FEB868ADBAEA88F3785C000AB22FD259A28B27896587CBEC6A4984ABB2D94E3F65701EFD349A64762E37E854A674EDAA7E7CE769FC87EB9E32D93DA0E42BF8745CB6E39BDE78950A116CB883074E3A97802952A838A34D652B4B3905347BFD47023EF2BCAA7E5C7DE88EC317D13610D85433260BB41B87A2A9F87D327AC5F45434CD3B58B6121BC448D236FEA2F6169FA5839A7475CFFE8025A32C8DC303C72790F24295BA4E5635062901513FFE6A21D2F48B94C5F3CDC3761E57D136E165DB0BAFC8E2556C96929DD6488804903E69A91261FECBF7A84F24534EBD31615FBD1C50AE3199F4935CD4FAE67C631EAE0951B0B7984227E3A4A05751E26B8A293236DBA673DE7F21CD53AE2719749AD3F9078287EB4F3FE3462ABE4F42D073EB7612EFB022B7256688AC05349BD3F2EB33E16218C156DB34C5AB4E5B0D7D300C8E5AA1EE012846EDC615A99C956F44E67ED270A60A51D298483B287B0BA3ABDA8D94AB7F93F355A260BEDDA5D8CA72D763F8D0B4E99312E1754D50D42A6CA1AC9D4A856E9186ADA36964D9E919C99255FEF36025AB63CF182AAB8BD4D6C8DA30392186621955EFAA03EA58834CCE04BFA33FCBE3CA6B031D0D4E5096711B2BE780A9851120EE17BA902683140C3377771C1CBF7DC2CDE8DEF3FECA4FABBF2F64462B40510B99F2924FEAFD55D70981D38FA983F86EBC5B04FEFB80DCC8466DF9840CE86371F100CA18388AE41812A72A34D9F886418C969BD96EE3922E5A56C37D3168B578308E5B62B0CCD91CE1F998F1698596B86317F78FBDAB601559C86709936B610FE0EE0008B40B1A51F90898FAEAD02550101886E953F7A4590A81FA08F8CC4A2263A0551088B8CC395BC3AFABBB702280172F07F6CB5334FF181F06CE15AF908A3E55DD0ED3985AE2591E8DEAE560CB820EA054927A1F79275C58A577884E4DFBF42A02BD5752B30A2FDA5884A962D8C81AA91AD955444BD013B76866771F738F047AA5953E3A63A740A065C06951EDEA03F34AAB2B878B8D63ABBF96FB80E434D65F8989502F206608EA95B6DD8974A8A31DE8073B4F4FD3B332116E8CAB7B30B180560DB719BE1DB825428F3F4DE9FADC12A13517028FA315EBAE4EFF56F195B621EC6114C2E635EABD5331AC63F329AAEBD5D26AF3D3FF4CE519CF8EDD848061C3E16E68459A99E9DD4AD5E583C47660243D90CAAA06BEC0E29D29E5DD02BD1F346668C7E44DFE0D234E6B2B85682A361B514C0971CD34DA844AC979E52F2186CB3810AC89D9389F4C52B7088188CC14A6559C7E073DC4DC2FBBE4A52692D6070EA821F82B65EF7DB2C1AC3830C23D7354F68CE2C472C3A1AF710029A2D4C03BED07272A5A850F3B7314EB7273B54693125EFEED5B16937460BA41EC74A9FCD7483F36D949C342E146C285C347D65CFB91D6E36B27A5D88376B89986A5327360B91F4972C24299C4301B26FA960BBE0BAF0DDACE54E525479C2331A426972AB6BDB5B5D1AFA5E77FC7C059E59E8D0428846A459B8BE147437AB721DBC06476B1D9806A4031BA3CE8B570AF0FC150385EF53C1FB257AC758B372662E92F1B2495DC1E912CFBE039C986FD9B48B929EDF601774CC303918BA46114899A4E29BD0C6F0B15ECE5FA86B3AD3997FEAC2C6B124F41FFD14029494E2305B71E8F9B8799D93DC4A0242211070D2D0D5D4C78B21AFDAD6A88AF72F500D8EA4F13AF8839419218613196D58C30979CEAF625922356FAE681A1944FEC2EE5D28220BAE72B01F0042E2521819963E33FD7247F3766031CB0E47DD052D7EE6F8A731D0B150F02FE414F314CBEB849EA8176710311E91A88D15D1C301A8188EA2CE57B23B30661BB9DE648BF55855427A0DAD010E833C9DEBE37F6D9521EB1493723AE951FD5C74C2E6168B438D7550F93C2C33753A9428F594330D9732C02678EF1095711355FFED0F6790A3F2826D1A003D926F94356A0B2B33710FC21DFC67C9326362E111ABF713C14C80E826BD864649E1B5258FD3892A35CA44F19FD287B0B0A3D79DC88E0AE5B5937A48AF77624B4A632C572F70492A534EC39CC3076430E060753D111C1275243A304E83E0DA481CED8FAF40B22EB842563256C39D0F2DBAFCF50B521625725DF26F03166FA44367421A0CDC6F541933E86C32FA1FBDD4339EB971DCE9DB6BA360E1EBFCAFF6510B35A5EFB67334227F19162C125F7CE805ACF024C7D8C295C4EFBF626C230F203AB22FD1DF6D4105528B82660ABB011CB334B626F292E05BD55CC37BB3CEAB1D0B32BD79A1CF3F63318408659FA4C6FD18B014685ABF43055BBBD8A70EF4EAD56A22E08AA1860AF5FFE1EC63CD83DD2F6D678BE933AA605568D0018C6F930F4E16C34E8185250D96D2D7261048BA5A77C03630BB1B6592D5A5632914165B29A248CFBF0EC05CC71AB9051F22F87C435457A9A1CD628732892FC46C23296901E4B831BACDEC6E35E686E485B650E5B5F70C3973FB944D17B921F382B8A987953061C7A4F6D740E6DF96C3D06BC046CDC872098CDD0259C0656244F0A4B4D2ABDA2CCABA450452C743D6EFAB053ADD3887E1F09ECF188F5BE39647143E2D7A4DF7B4BF03414195D51BEAF5E8E4EFED3705E03A2E55AE4F8F4AEF920A28048FB1D27C91A5ADDE0A457C43C2989B124DE28166551FFC64AFA369694CEE5088395B61D5CBA1C151622843EB1DC6182336539E86D6D8777A23A4ADBB3F583F9A309C623E0AB337CB184B9226AF845F1A1A9663583C521FD0554E86B49CBC39FBA8664EA6462A7F17D79061BCFFFDEFFD414AD51C9AF7E0A8D07FBC15142A96A47E071E921AC7FAD475E884617BB38BDF0F5C0914B2717F5B73E14275E1B8278AD531E9E17AB77C18C2F99EAFF50F54C7DA49B60FF1BBC707266582F2D73C7AEC4E6359B115D66DD51F69D98DAAD04A6B8215DDFA3B52BD2A5AB18D8852E776789EF48107954746761E79415CF7712A2FE16293DA7DB6FC2002FD66990205942332AE40645FC5465A46B93C29D532C7A971E14F9CB2AC5F5AF09883377C4097A24494906BA371F37B2B79F4B984ADC79F2B8E048B2FAA5DA1B1C67976623425F50EBEAF265824FDC06D40B192C9ECCFB84C449B46AB12193912438FA9C81DE66752EBE93990C3AD18CED7CFAA3F104C0B437B855C12948887B500C1A3249C847808E5835AF81F2DEB61096A46C13EBE7CC751063F717F77688F15A446B5CD42CEB3D5F6B3BEE423164371CA629EA70F10C4BB8D34C0C7B96A012E52F8367AA13BEA86A6F17C804772E23CE9D59026D62B12B8B685583F0B75F6511561B697DCDF173D4496DBAAFEA304168A317F6CD2F226641778FB9E0040DE395AFAF4B5638388E1E00D9B72EA0A7DA94012FCAC576CAEB9D72A2AB8B21F31137F5E44E8A320B8E39BD5FCF124CD358A785B93B9F438776DE320D65D10CAFE6A31EFD015C01E8D025A98EE2DCC5F642533E0BD0130BA37A67468753097244C374C0960931D7FF2B166E3E3D1BB6367A251BA4853AEAAAF81C9715F76E1E6CEE92612C8E4BCEA77BB83D27C1F1EA56E2349E68F6C119FCC73EA53C60A4DBEF2792E43DECFDEF196112B63A71599F20D6F3B640C377FB11CC385EAC7D0030CFB3F05650CC447B97EA46CA4A6742393DB4C067B8B100D2646387215442FC30A435116CC4246883711E1FFFA692B53DC13974FBB483C0037ADED4A539231D1D6A79F1CA7275E642EEBF7944ECD7E9DEAFA53E4BD7CD88EE838B9DC67238BC1FEEA9ED8A45C38A52C4D732AE1D9E6A44859867E0C6298C2626DF7360AC503AF49030C617A0ECB29183AD0618142487D7B86C0BC92595D58B01D152996E28328B3ADDE903773757F5345EA896F84A6AB843E61984B58F1CA4F5F387A8E6FA7896D2B222C326935730CB31FF36E64C4DDA9469DE46FB52A2C1A26CAFF005A7C33ED2E9377CAE934A6C41C2C056E73C6141C78B4A0524AE3EB67FEE322F93CD29759DAACF5AF4D8763C2288A75DE0FF1C7138D046FB37A8FAF98012C4D0A6CF3F4F0D3C531AC428EF27AED0C269F5B77A4AFA58EB94EEE68D55B0E27125A144C71DBCD940F0FE6E52189C1F6DFA051DED12714496F501F4543E788735AA0331B6078AE9D6E8224B3F45AF639006FB86B393CA3D529F1F326E446592E9C91676013A0E29F3229B4296168ED77BAAF87B0A2BC63D5844587095660329E0F71F12ED6A17D0DF6E08EBE57496D385D14044792F421AFEE5E34EF62B9D37151A6E15C99A1482CCC14B91951A041CC655ACC662066FC53457813FCDF5FED92D7543272064A8FCD71ED1EDE472D140010538F27E3B9E51F23928D16854F6907D392B32C48C6B4B061FDA6F0D3AF16C9AA20B054A309D14BF45BAACFB18EA59BBD067BDD8AC6EB7474FD2E4CC9059429B291D4182C7A6E38FE9B2187C1A21F601A0EB63690D7436BE04DD7418576C65BD8486EDEB7FB09C20BB417724E998886F653FC2012956E0618295DF85FF069B26432331A9B71E442ACC4DC6327716B4E414D1F9CBB25738B3E4B6B74DCAB67DA8CBEB1B7391C449DEE05502853D96035CC0632290DDA2BF846D630E7C0F630AFFAB22F924880AC3C87F1C1111D744087D507C1709EAF0F0A0109DCF92D5B90314B1DFB51CDA2410195A2C33C22A0B252A9837291F3735B3417689614A51ADD81067C3E4A712B1A75B40755BCF3CDF71634A8A8FB102C23A20E7F694C783E5D8734ED3764CE7860AF2EB9A10FC8FEAAE7BEAA7B54EB9CB21A27424660A2782BEB7008C5B873B6B8928F5B3A91EE253A5AB58201AAC414043ACB70EF28964C323D8A572B6431895869E0AF7196AC31C2563E282E36CBC0CA39C091D48E57F77B2F8813FCF8C0E0830279E30394E6809AF95BE8DA6DD3EB3093C60AD7347F4A5EBE0D423B46884FD48C20EFC839626D2F0CC412097987F0CA5DD16F5F309CEF0425FC839D62A34F86411D53B796FA232246BF47CFDEF71B973C0D353C38AD66BF19967C30112299BE8A8185C6E5ADD8F6E14AE30D53CFF766B364DF4D3C74E405AC832501DE9BB37DACACDBF1279C9ACE81A2286947DC023CD3FB823E65D3102D675D396071FEE286D34957744DDEA2063D1B096314F94C119CE88E65EF1B1BA91EB2C90C7A901DC53FD84320D971F08A5C1BE1E72972B6EBC0FE361895F602BA42320F5096E968CF8D3D097DD2378BCFB9228650A9362962579251A35ADA23304646072662C696803221010E5C9862D68AC42254EC74370F23D98BB14D0D602E8F81847305AAFD1C1381ABDF2EC08A74B6B77711B8797082F93AD8B4158643097A6DC9E90F819F499DD06229A2F187B6815ED9DB742293C1F5B20E942DB5E45D2CB54203FD0939C65006AC68087A0899658C6AC93BB604DB81FA0BF8E9BD5FB7E74F95A6FAD3883890B681F28AE157C04EC267574F84FFC713D667C39B41857F6572041868C63104FCFF1CFE4DECAF589D5C3072F5754113B760D8CC7122372508118625C9D11BBF2C958E45EA525B5AA1AC94B44892A96315CD72833CB60C88456B9DE2FF47D9DC5A726E40B55AC8E60C9B1627C749F1CF2D0DD72AED7C2510FABB637A8F330EF09B1C768DC73C425332A5F430613B7D3A3388A44E2163BB57CCA046E0E88F17E082F56D37EB652E5814D344A2799058CD74357CA24972DB96DC1C0D6B4F8CF550A1B536A05C4FCFFA5B764D1BAFA74EF780D579DB8D5B2F6C2261B232D3DBC5F7B0675C93BC29C4E332BD203BDD9D5DF386E631C6B93DA810246AD564358BD3B822B825D7051E3025E234379B7588BE86B7FEAE044BDF9EADD3371958AE559EB0620D7F4E61FFEFA9F0048B7637DC81E1EF6045473DCB584519DEEFAADDC32A0ABB66CCA5A446E327CE97F82A00793075D015ECBCB0D2EDA84E54717D0F097B85A4381F8185825238435CCCDB0A06371B5E47470315535A845DA2BE1904CA7F7AC59A2D057D0C12121AB64B7161D802152DECF1DA5DE4E222A49003528F24425A8DDFBC1E90D4FB739FE230CDB116DF7D6F4334C8C1FE8C7302745E2AD827BA7CD9F64B8DCC373DA80F6AF880387B908F8960580413C21375FCC90FF9615E683A117AD43814ABD5108C76C17C475B4A455EE9563EE4285A9421063FF28E05AC91F7BD106A3EE60D9D97E250944E691480ED60174421C1C45CF5DC0F81995618B1F03A08FFC0B1CDC1526AACA41215EE8862D23B7B85D29FEF8A6BCE29677C8BF17BFD857E99CB0E548E9FA4AA20481098626A3E0DB838259C7B109BFFBDB0A2B1FB59A3B329284BF7C34A89D0F5BA1BD8CC478C0BA0618E946B8013E36D6521DDE598F3A6FBECFA9CBC25368387B1DEE7D28AFB69DF0FFFD71DCF8841E41A995237ADB5992C922468073DA547174F2605D63F648D3617304360F8480265193D569B66AFD7F04D15BBCE8E8FA4F92C6DBDB693F7DD91F944D8464321E3A9CA0654D6892D37C5CA1EB671726374D3E176D05E204A1BE4FAD07F7BB0C9D25761D49694337EA3EDB03A294FC1E5D83800FE03663CBC310563C06F9DF45F5E5C67B7F5C1F766B7B4576B80685736C36A1368FAB2D23334DBFB9E20AB123BC8C59428889164D3F1E5ECEE0B2D4B7FB2F013648EFA16C60306D52C29859EC1985448D1E40DD21C6047A6DBE49BFC26936318AD63EB1D9F615A6DB5CFEEA4FF48B4144AF32BD60241374D697946F9E21FB3D7DBEAB6F1122070169C36408C9BABA3B5B2F4F407409AE2F5C238A300FB22F86E1CC6825BABFB534BBA45DEDF8CD09758A38403EEF292B6508152C11D6EF1F57E0813A9A80B19F691490B67AEA73D4260E0B4D0994F69C93B1D752861E69D934280E5E9D2DEA66ABBCBC03D5B222A15B58A5F61C853BCA885E84D4F72C5535ACF584C027918EC057D69C005F4E223FB4AAF57A3FDF9DB7E0D1564FAEF5B5CCB7E70E1F5F9FEC5F5F18FC4F7A02CFB8CD28FDABDA2C3FBAB99015BC3A5B417E7D740D605AAEAABC126B9E902CE4F9DF210C45D4A56F8C3A012B8AE2470F4DD344ABB8F09E7FEC6C8B9B4C85AB415680EA1AB6D1E8E150E9F4D1B8D3EF398B2F99C5F2E9CB2DC407C2D0062DC59309B6F7DFACF83C615D4F7AA2D4988A266F03BC1D3151FFF3BBEC433164619F30299491B6F537052EC199C99AC5C4F2F8C117B5497161E80A604EE7C7F7B29A124A984DAC51D59AA7E02F51E097824E4146F9535BC09B256E8710E5E1CD5798B96281C98F31FE4DC386017B30F42559DF13D508FE318E16CDBDD8C1096023E907B9875A27B9D7DB32163CD885157013DFFC6991663F6897B01A668D432218B6BA1DF34AC670863A963ADAB63E0A32F27E9EC6043EBAB4CBE872CA9A9E1BDD1D6EB07706D35894FE2C7BE905FEE0E767B1157E954DC5B8FFFF66BC7B558E4738D20082AB23A471F223D87B69548A2C0D23D40C0227EE1163FE0C2632D064448ADADD6CBCBCA63DDECD7B914312D03998DBD1144EF37EB2C10AFA268E9BA7495CC28048103614EF46EAD888B805AAABE4D512F821BB8404253B379FFFA536A45576B25C8E5EFD228FB2215DE54817F62479DC4F4E8E98960275D65FCB8DF4A5E87BA65BB45A6781B777C324E5B5D353242DB288E6CB738E1992776EB557582E06637BF603543D27B27CBA11BEF936C6BA9590636DADEA348EEC79FD151262355A72E784DDE81C2B478C417CB930B3A6469E3C3C44A6EED2045354C744F445B6D4A2E80BCA0CA49F40DFBCFDC7539F111944EF46C8CA9768A552814FC22AAE28D9E123342A9E52EAF977DB8E76F176A697EFDF94B4B1050CDF26B4BAB1C64A3D11542F679801ACF24867A403A007158DB3662BB46149A8BDB99B350F4ABB1BCB85C81C146BE25E684C18BA2FAF53A0E752B1548676BA7C0EBEC841E47E70DACC127E185C19142016483CDE75E596B66F5F58549FC659FD8C19A6079880B192F33A15B88A0714A24B4A92A9AE6F1F44E734271FB964FEE55AF5E65FECB97740D57DB5103829C366A50A2030E1B1841BF0B88E43635AA9961899C1DF8BF032EF6418A1E93F1F161B56A94BD08AB81B36614EF10A515057498361EBF8686E6409407AC5AFAB03E16D365E9671BEDFF6288F1AF9BBD907CE6D30878EBCB906209227A237363B3B185C98C7B4308CAD3FCFD525FA6ACC8D7A746309C56F9447E9D927D04B36A33A60B663C005810E9F07B2EF9ADA4A5DDC62E2E11C4CA2351A1F21694B8779F9B59EE2372D5C6F1E865CEC5871F830EF2D001E37D2C86C7B8DF874500D877AF6921AEB0E4A1F021BD7F78BC17817D8F4F5A87768AFDD0532BC7951969F70D465F30313FD2D253A4C93874051612B7D72FB938FF6736DB323B7349ABA23E6538B7273937E0E8E96826C5D8DB9355A0DCFA8FF790F3C14F5040511A4B94AF1CB242E46E0AD600EC187AAF27F946CD1AFEAC7342E11D9B1E24CA059F2A38378309CCE69E1D673FC9EE2A32D1682D8BE580924EE8A9A273C77F165E6673870A47DA69E59877FC269312461320360481AA4E539130EA12294BF66320D38E48737F8F96D00A29C162ED2FF0623BB60566782528D2DAAE912C79F7A15CCCE0EAD05C9FD0968EFED15979F7D67191C7CADFC9CC954AB75352E4794A030FD4604008D6D15EBCF24D5ECCD514541697643E7F975D22F8821F1DDDD6AA5C6587B1C34DF6E78C5AD75F57C703AF6A689D029A78ACC74CBC9CC25A3D631C60985E2C4BDA0E8A0967FA464DAC3A57164BE7346187AF2654DAE213F7E8F92128278C9C9838B66EE30BC70055B3AFA9D69FD103EA6516D67403CE96BEEB727EB734331716C65C95718B4371E089F27E14676D497F6064F3DAD6EDDA587F22455A92BC914C0F03A120E1286220DF3F4568F9A32B54FC1DD203F97725BB50C38D49C7B11F29D23912DD9CD932F710941667CB03DBC024FA7B1FC34C875C8B8FE2E01042F37739202F998B8087D5A10CE3D0812D504CA8B4CF249C1D593DFF3CAD4D58EFAE235D33A75E2EFEB8665384BAF3FE544F7950C2B8540CFBEFC4F89B5C14A478A6A0F69F757A1AE1ADCF8DCA3996BD58E3BA9618F6FCA558FDD2019FE549339AB3F740F21619B9AFEA8D7AE125292477144630427E422B5C72EA721F84CA889F817238F088447922662995ACA84F210319E8BE0448639860BF8BC78362470AE115EAF966CD78E200FD0F5672D92AC8D886BEBFCCBA24A196DE5326EAF53719558B870CDF2DD8490412095C7A7118E6E15658AF6FF38B1FC2F00E6FEFDC48CC58C62739BE65423EE76E4239AFA140EC9B3E756F7497EE81309E5D08A1556A8D1B7F6CEAA7489D560F4362D7E5E85FF84FE9B6293C6D948F1D603ACB27956FF64019FD3381B582E8F44C11F1ACEEC86E9FCF09D5C019D46AA788595F8EF0D58220609D5F6B9228CE02DF178D53BB578DA947CCAE428259F7F1C0BED436D798669E7DB31E1B3FE175464FC671047D2B178249B4EF259149D5C8BFA02183198CA586FEEB5EB4DCB894F16BB0A3396EB12897D2A5E97D280F8B5F7846017AD002FBE261D7AB2DEBEDB7CF569857278959DBA5F20B4BBFD7944B06DE4A78771F36FBA9F0FEFB05DCE0F633A174B5FD6C152E5753D6D3873FC7DFF41D01F6EF69FDB04D8049E0C8CFE08929D9ACBC2328376E11EF06CB0D5D027948A3ADF22200952715F9C3702468B16D4AEBD9515495E59D13972B52B2FE724420085CE8321B540D4AFD1A5609D2CCC80AF2E9C3853C1DD1A9BD67B4972BD1B2170B459726ADD35A0B5538785DA85BB65FF20E6A7798E7B1B0CD9AA7921A4669D84273CFC33C6743EF3DA9229049FF841A37F733F792BF415F9FADA5E46D95F92604941140E9EFCD22BF68C315640FF2281EEA6AAA0779E1B110293BD59A6B0EA4B3E6D2661B977B9EF253877FAE03CC68B1C90B6C1C4297B320D4842C4D61852409B28DCB5D491397D5CCDA14AD7E5ECAE440DECDABBF87D4E1C5EBCB059AF6E7E3E5FED0B94EFF3C374EE885DD2028D4823C18636075395EB4F89BE8B5E060EB178AD9CB191B6AD68D79674E0101B47CEFC3FDAE089CB195C53D75043BADA6877AEDC5BBDFE1E863272F8C4FD726548AA989A65FBEC9463F8B5482CC75ECE46F7260AEF2534015EE82633627458D4C263C8CCE27DF97ED39288375D1780BF46DD0E7287D02A529AF1568C4408D6B8C82E772ED99CAF55BA2C9FBF27EBB8DBCF7F270011E1E76E59A7696C488099CF1FF8107CBD1DBAA80493C7932CD64D2A17AE84E897795906739EF47F6E3C57945FA8F6DB1FE9233DFA3265ACBDE8703E65A2A2DD550A5F09752733FFCEF390B292A7391342639744F885309A78F66882B6EC106898558090F463A23928D7FE5072A13408ECF5B1B4B06FEE10B6E7F1208C2F307C412FDDB33D83DDC6838D39071EE4FE8D8AAAC82563379CBA198FBF03E79D6D1B1E27F7A15BAE729F336023C446C6179223042A9A458A581534319BA181993DDCF1D5F985F8E9A4B92E99E8C9B4CC7E07EF098650AECF7A7861EE9A5EC172E066463552BC38CEB3EE8555770F6E20F17FBA4FC857B54717CA33A12D87266D5C818DF95FE5D46413B51831B4D1E8587D53DCA16B7C85ECA11BB95159609DD13B0B68AF51679731D5563820D8ED2C15B8CC3E67FE596548CB00794FB7EC342FA3F4CB7F42B8660448BB05F32D44EBB59184967A451EB817EFC4698356FF073CCB94E026397EFAF7DDDD40CB6BD8A2972158C60344346F73662A7452A5C1805F10EEB45E02375CA986F43F6FDB0473A7EB1E8376B32F2EF2282AD2D0E60C1F2D9D55F1B5882BFA5D7CCCF030268ACEB3DD746B3E287EFCF105554207A3495AF8274B189CE2161DAC99B66D5887596DE3EB8F6BA50A3BDE4ADE5FE23C6AF93DCCF53F0927527E21E1B449EAEF31EB3A3BFE2F821C210256D9E0B8D0353A9D20DE2A902D379CC4C90E2590D6F2626416788EC50FB5D55FB27FD1C96765D528386BA0B101BF1A74950C043CAE16FD167671AC9DE31D746129377604D2CA0A9ADBDE20EA8FFF6D65D545269C708879DD146CB6F939FA75413DD732612D5F9FBBA169AF7F076D94E4EFF72D0D95A1EC0A1E1DA34FEAD3163EE229204799290B9DB9A6B250F23037C5DBD1ED19E0CBFE26F27B3BD7E62AA214DD3573BB54481EA7F5F1F0333456DE9071B1B1545456E6930CA281D5F3815EC5193D73D98D328BA35B14DB64805D51DBB77C85E59266B457A9F4E33B85DD78A818B9E54AB6E44A29530AC1C648566A8C3F24EBFC23AA46A5A982E55D9373980AC41917E28DA236DBB6D8AF77D728843C815584D750A3740BF1DABD3C70CFBC4F617D4283111A203078F50AEB966D0FCDFEF92842FFE8F1A783DBC90A6000399B6929060A9E7FFE28B65D1E86B0CED7B88B7A5FDF5760882E181F2E6AC815CD7C3AD64F09FCD7C87D9E5FA6C256782AA2FBC953E106C7583A334B74DD6C79D3FAEE343C9D44C47389A5991289D93912EEE1E121479B933B5520795F9F696CF9D245A332DE5517A8DA46E04B3FF63D97578041A54B9C46CA468DEEFEB41059891A4740C3DCEA0C172AB97BD9DA2563E44FAF1CB59FA36F01CABA7691EE57228D8CB5A25337E93373D0F1AD69380D76A286ABA63891958EB90FE0E639B9C713BE8D545FF5570543F99A16E170254C737DE2553271386E30CF350C6769DC316C893559528A903BA983DC4531E52A00816A73FE5C3AB08E6509958B6B9AAEDA1939FA1E9DB75875044C867364B583BE35A7C1341A0F3FBD468D8888128467A5FEF281A1EDF3DEB7CA65868223D494083DEEC2BBCF46B22B68652C06201AD637A6B797D8CD5844909506C14441D52DD89D291E3C82A748B41AD2055CA244B6A39B317BDE06AE62918489DB31FC1A1805329EBFA3B30135A89037A512FA8E8E39BED31F45ED184BFC89E9ED340B1E6ED5FA327620226B9A02BA89D4DD3F209083FD6934B816AB7165834940C0ABD688022F72DA8C09801617B800BF5C17F6644C5905307811CA759C61793955516FC9482EEAFFD1029953E77A42AC50F88E1448CEF013E7DAE4D02B45AEC084F953DEC1305E0FF9CB87E39472BBF5B7E59E19F22114982C3E33DD0731C1E592EFF437ABC37C7745AE2AFD3D725C98713A6697CF054AB135143D7B142C5BD03A52A8C0D76C73789C1638DAA4E9E33FE8A04CC9A73112D7C5B59B535F91A7519F8207C13F6F21A104BD49B906A6B93B28CFC41189F0BFD43BB357C6FA923B6BC06608C1349AF70187C93ACC69F6089C60EFE51D3677329A1E32C63A72FF1EFE50B93931E6A823D092ADFF5340B33C31AFBE8A0DB184EA7D9FFD6FA488AC62F7F21D8A4579470EC6DA52078F8C79B56E02D488654DB0ADD6C4D73D7217364376138795E470FE03C1F163C5068D2D8DE065E0BBFE1D9DC5C9D5751BAD2FF7868EA926A22E118EFED6DACA37D81BD342594353CED3AD7D01AE45243BFE9AA32ECD14EC8F66598E6918B4B133DB894F137253A980C57D3186D652DF80D979FCF582407BDF72A100380A56B009F2E754F29CD77A32920E999C147E315FB0DD416A0146ADFE8891AEDAEC7FB1EA59DFED3D1C7F30F24D7D6A9096E23CAD39E9C889B4448BE7520C76389BDE7D6FF096B58618E5D6CE53B845F1EDD6BA3A6E0A0BDE6FE44D72BDF7B8AFB27B71E42C63327BD2E7C2D47989256C037B3E1961B2EAF99461EB3115423103EAE6BC104031DF27401E399A0873BBC2B5B3D666A4325C7CDFF088DF5CCFC5F5F3CB8EE26DFDCE14DA9C0605B580DFA5EE47F6EDAFBA53C952F0A9B31B30D98B7E963E502D6E1809410E349C11A23CDBB053ACC61AC86BC8607C169B1CA721B982603BE98260BF05E59FE49BE0C84114D1B4B56C39C9940950BB464980486C3C82F210DEABF8D783171F91DAF78D70788F7D945AC2435317065B0285EBA65289D88C98AB7CEFC5103A87BF577E9ACF133CC87BD9F6DEC3A82CEBC4622337A3062D0280EBE5C50600D6F66F305A92082281B88F26F302BAB45EF2800F2073F8BEE2F2BBAA3F45249DF003D97ECEF16993E91926A80CB9E7EBEE44AEAD876D8DD49B33A40AC0CD6C1B628352559B71BF21950E014BB7C750FD9DEB2DF6D559B86133B6344428C6D885415010EA4CEAA0487CF18A77D32BC6BE9B8571EE233ABF90E4830958AE34FC30CD02F8194D8DC3241F051331AEAF1ED748CAF775F47CC81A8406ADE208FC42EB63268DCA948617F83C4BFCC51AA178CD832E303E2FF2947B7B20BD45D810A51DF2DEB14CEEE39EDA0B432D369723D04675CAC41DD77DFB1B4CD77A5E89FEBC171D664D581685FDA29B8A7284D22855284AAA2A7ED4774ECD2867351B9D2DA7FA7B6F364CC91BBB75B1F1035D12E2AD99D93F4C527CCB49F43459A417F46CF8018429E7C0550947223C6260E2355B1B19CB9DC385A4378D7E4EB19A014E04634AFA3184C2E39C05F04A69680A1C8807555CA4F48008B15B81A98CB1EE08E5D190E8F0C7FDB669365466FDAECF1B1E46B2B88A41E5EA7F976858561A711B494D7013DF9434630D161B4EBE3376CD672DD9EBD18045969A2A1F5FBC79CEC8F097A35C74003B46EEBC9A2EA174B6C07A854551C0314E240A3629505048A2954FA50CF520CE14C65607E014DBD7F450461F5E0A685534B0106D83EFF119BC5DFE7CB77A0518E85246DE8EECC1A26B3EAD71211DA94F72C7EEA8D09976A583578BEC3318AD44C0E4AAC1E8D6C3F511243C8EFFE9866265810367E7B74A0B26A269A3692F76D3D58622B47185C2E59CC8CF0BC6E2BB23F5D80000D033AE6DE3BEECAC16CB253CC8D5A45DC103603B4849F82E85E0E82551566E872A8F5A17B8E8C13C13254BE968E43DAA5B80CE7C6A55CFE74154FA35D9832024F2400BE24F10DA65CE4E71469966F311F64E9A8EED365F5821299BE64F491EFB9D6247730A7AFD0F2C45D94F3C58B5B17F1359989392EB9667A53A34940317B408D68FA3DF22A40C4BAC3A0F4EEA159A4B0192F9C46AB2FA0CFC4117AF4EABC2B766DD5BD01FDE35E2F0E2DF5891897E01135B1B07E778CB407CA2C34777FF2D1CD8613A70DF02A81B507721A02F118A2D19C795E65EFA4542E622FCEF261E927C75E48224B6795892A2BC805EEC895CEBCC5799DE51CA4E25C41CADA71FB0886BF47F9F4C88CC3A6EFCC7B25DA00788BDCBFCFC3804EAAB76129E3C1BF20D4A81D3B3CC9AB780E578654DEFBE03945DE39072906CAAEC6BD7E190A20E6A9DEAFDCA2A3D54F333DCDC6B7F772E1CDC0CF9236CB4E636B5F84A081EC5489D675B2A2A0BF874E52021B6EDB973DC9EBCC194F28F72A6854C5ABDDB833B9B593CBC90B8A9038F0C5033495B62A3906AA0E9C06EA6DC1AB4ADECA8BDAB437CE5E263AB614241FE35C9EA7B4C5B3B7BD6A96A341206527F6D76EEFB9A57C364E0363DF76CEA10A09502624A22CCDE4B50D3AB3AEE435F88261FC393767B7BE9FCBF4206554A9462EC2F298B2691E3147DF3915D77B2D9FC5ECD54C763DDCADE855BD7E4E2A2AD6CA62E7C5D798B3760598F2974C2F2F8C4EB4B3F8CC71138C336CB433DB9D4B90907392E3B83C5B0C375286D0231D98904120180812BCD18781FC25840610BCCA4FC8640A5E619B4F8C79546BB0E0686625B11AB2868283C103C00A2A9DA1C928D5BC3DA89E451D5B742AEF201176388CCEA784ABDDE6342F6456D578FD432A068BA90EF0A725A457E8B43AAD56A9D2586E16829D407A5F9A38E228785BB946AAC9027AB4FEE3046FD96DFC7343A077B8CBAA47ED227C45A0F4025C00BEB99F545499DAEBADE8BA010E12AC3F5506D9F585F2EDD2747E7EE2AC65FDCC188F936BB7E397C85EF880AE8DC23D5BB63C20BB917E4C1C6D024AA2B2DC1847EC9483FA3674B3F9F69D60ACB4F38D90EAB57729A7E015C753C14EDE909B3FEF9E6839C4F7720EB15073C8BDA7384792184B30E1C0B0C61C30A68FFFADE1B5618967C5E0FF0B113A14A536F491796DDCC641A3C69C6DA76F6A085CDB001B31BFB469A760E5C1BD3F11B3B9983F96EA38A79A9A1E724EF92E06C844035DF97FE6CA600AAA4061DE3641BDA2B191F6CBC5500ADA6CA9B7A7B5D00E1AC17AB3A8ED71CEDF8DC3AB978FBD023100E07BE8E764EEC0A05AD335B49C57D95240CA2E9C5EBE960F5B1086EB6B9EE23EAF2F3F2038B68717787025B133C7D1FE17AECB5E04846F61792D4C2AEF45FB5D7B0A67CEF1543A02AF056EDC270D7D6AF517923343DF4F9BB86978E26F2DBA8AA8F7CF97DA3646E9CE2F1B9EC0C927BEFB35904B7D4652A7D7E5894E8B0C54BA6B3D9C717C2707C16E7C5E4B86B48D0C9EF654F1422E062D34AA6B362DF23B96FCEDC0A48836CFFCFFCB3C2031C9885BC893AB9B7F79289CFE69AB4396A39D2CF7701B4C3882D2D74928E2FC9F2686666C874B83D24453F2CF7F0C8A0D63EE8479EDFFF5949E1EE00E953CADBB992394B1286D1878FF8DAF6EFF1483B8038C65D5346FF0266D25D0F88245C7E1EE44CFFD3F8E359D9E2BB60A3C8FC353BD24D9AA25039C402B9BEB98E17066CA509AB72FA04823D5B27B568986B3F6C01A612E44BB1DAE38A76D64F2C28A8D18C715DB3991FA41E369F3CA392B26CA12A8127B3F78D5AA08BBB2F3B4F5B436CC1728BFFBF23DFC8BEE255369FC241A6B67DA31E755ACCDBA279BD0F1E6F9226A066940C855551B5BF4924A091ED2A1206A4178DD5C7B79710265BA5FB300DFD96394D15F07AFC2A4352B50F51F2C593D098434E2CE12844AE2C33D6B2330D1A789D5183707C951D878E8DDB684B435703DD8BBAC3EB692766600EE18A04E9532CF24D4E28CE2D00EADF172F7731C7CE2D1F9320E77442B6EF97CBBBFFEC947B3791B40693B3E722211DF9FA3D8C81AF4389EE63C718293965C825E37EC8B02AB2C238C5E6352C8F953CA0B12D09E9643F2DC384B5595EC3E02C55A97C3F97E5C989B3561634A11623D84686B75D8852B7F1759AFFA89741CFD64856C880CB7665B123BA902BA1CCBA5FDD832645A47A0BDFF24E7122423987F9F9C7E65D2C981850DFDD4C928DB466A800594695F80B1E1C64CC4918377194AF24E4A1EEDF3EA85EF534DB004E621D65806E7E852B447B0B63BD96E602993A320D79FA86754E32D36FE5CE8E83B0A446C56E56F72EE7E5511630A759D1B089CC0F9E80E1059AB28F674025A8C46D784F87A2298FF799E976440B723E3556FEA98FE838E9F8093A4FE668B59932CE569AB30DB4099CCFF49091FF16FD0AD4828C431B35CF59F87C29A55D955355035C5A988A99A0C4062254C92BE0DB46B9FB4CD95D345074F11D8CBFB7E6D8EE338F9393B2F63EAB0D6C7A257CD1BA5906B8215D88234D7AE8C22069089FDF31546AA3F05F81B46A59D92804076608F43F64C52AA2E6EA2B133398F0A2E3FD4C73D2C716823C3AD019C274B2EBCBEBB7DA917D72F5C0E81AAD30ACE3B0F8D3D60C46D3AA96B8B3DC662816D56996B676C82EB182891D1124D5C67F02A0408B3C4043F9550A8573D11ECECA126B47E143E7399160427F19FB30F61D50516CAE025E2C360E9B5769E7A73F3879021E50769D376DBC4A97F17E5619A12E1AF97DDE035FE657E9F130239AF362089AA48B73EF0B7EFFEE32B03E1BD8B0B8C8106FC6DD55C3F3DD46C714CA5D9FBE8A48B777015497821BB733A555CAD1DE42E99265D0AD849EFDF48DFCEE5988E1868B523645DE1D73775EB611F52527A123659D3D28D8D475A33FDB50E73A52A46AFDF51DFA415BC452A8C03C26F474EDCB19A629A2CA8307D18D09EC1F2007B1E881855075F6655E7F51366BC70D7F320D8B0AEB271ED31862136095979A0EC58850FF0B15E175F75A42C5F2282EDF523522C325C38810F848F1E0112A0F50F15E00A32D7B52E506E4A8C195C5A3FAF34E5F7127F128A55D62626AAF8C3B4F569B092B000E7D591C23EDD7908CCF7945233E96531646B49F1C9D8450C9075B9D901CD6CA38BAC85662780754F966119D97720C1A4CD6F1945A03183E11A9C4E28626953F0FC1A7620ABAB73186084A9D761BC8B1732F6723ABD0DE27DD52D4C5F074DE0F77E6149C217ED48402F6E2B4C824B9478F4AA8BB29FF6A82AE7FBB3D7369245E1FD48BEFC2B47E9E772F77DFC0CAF61E5620FDDBB2D708370D3FB34D497738FACB04558AA98E5D0EB9707774432381D6F5564845DFBE74C55157E7C591DCB82D48667BAB2497D73512ED7B2308DECC188252FB801B13A817F3B08C51E5EAA51179F45535CE73AE7CD2F3EB986EFDB0035DF978A814284C7DB814621D7AD14D2CD8A883E7C0CC57522F709F8B3D4DE2D0239995AEC44868CF18F545D348CD85D30ADBF2E6E2E5364D379AC86040B7E9A87D210D2D9FBB542B96216314D380F45265902C73FC7585CB893C4BE2A86228FF691436509B7484239F7BE3ED696251BD6F6DA3E5D8AD19A76F4AD1897355EA4802D1F009ADB1D7CA9444B79BC1A71D4497121AEF97AB5ED31BC9804222BE0196D3F93C6E47AD786E41B1D0AD95698028EEB8E69AA0ACC9B3C18B433D74701B3A6268B2FD3C9E9E1D7EFAF71A76ADA06201D66C5DA76AE2A4E6EAD4669733BFC6A5CE2A0F606EB02CDFE7B885BB947D781853C04F908795BFFEC2DCB760248D3BA29768E9A2B484454F905CA0FFFACC35459724331F1CCD55ACD786D879D812339D9262C5DB1CE8FFAAA9A4EEA2D36E4FEF7C556EA30941137FBF3197B9E5277184029884E47D335455BBD642E67F9500D4A3658476E5C4F67679FE98B86A212D2E0845766D923625C68FA231AF2F2E7E5F7153EE56A93EEE10E9F4A90E180F2A4295C1555758FDB7F56EC5F604A08482F81E17BAF140C345AF5AF153991D2175323B99F02D98D0EBE2F08AC231C0D58124DB1C046DF89666DB1933A7DCE86137D8287105607E325488FB1F18DC9E72D2BF642B6A613BD8AE0D0FD3364DBEA4CABC352C2DCD29EF496EE2688CBFB06FFF2F39F53828324E05FD9A830775097ECEDA4B09EF0BBB9A6DE5D9C7E9904A6F43C9B2C3E2211EC0131C87167AC92006D183F6E546AE425FDE5A57AEA5736AA493DA199537B2AF36372E6087AA1A9C906E33AF9E33CF7410C4BD4CB973F853005BFCC3FE6DD75D402E7CC7399A26D2B4D307E996D87EA24A1AEC95CD247425EB4CD5215857F85923E94CAF0B100443D194D32AA4DBABD3CDD97BB5FE41A34226D3B667CCA0FDA41EF8B1E27A074981B0E76CED58863A20905401D2AC71BCCF8FC6221CFA2F011B7EF64E085836B185304EA31DB1C31DADA384A98558DB146F11C0F6C6E2D8FE7171647978D3FFCBC697E88E8D42CB547E3F312D61274487F536A7F69CF070115755C91A251374E33B1FA37A88D8FF03D1D29260F169E9FD5B11BB0D6CCE10C426F87854F851DB533E3E8F1CAF50BD18B0E7C22145407350C6A76FC272F8848E5D68088059313288D880899A4962B5EA29E83BB3CBE5FB2C4ACABFB7F43947E092226C13AD66B2CE4431CDCB5466CCF82DAEAD6685F26E9A5B6F070823A7199CFFDCEB8541ABA4AE1F75BB67F577E9110FBCCDFC913991E60119911204FD7BF881D8F60555888B71FB60B19B07B8E9D1AEEA90725EF55B119CD1BC3FA7A94C17F1905CA874B68917F429D453F05F3956506BF53C08880133C752E47F910C5AA87BDCC6ED561D8C4A28A954FD51F8EE641FEC4521E4E11487B80E78DD4DA06685B20D800F9C701149571F63512750AAC60D7E9F9909F60A199600F255BFD9A5E53F6EFE0B87F8B706BC63A77A48CC71B4677C98CAA27424EEB19C6B07D84FD04269D62CFA349FF813BD398EDF606820528AC92AD80DB85A83AF00E7A351FF6AA1CE94A887A0369F4AF09CAF7F38D2D46CE9C25F8136D21CA43E529D2E15B5B56D550EABC29776570743E545A46D1D6473F6E43F41922AFB30023A1066C6F271F4575F19809A7AE571903FA0527A169C345BAA6D7639CF24889025E6042E7123081AAB1B49CBE85147D91613AA03D9BD5DDA3270247A8346BC877B927C1B07A301DD2BEF5E1E40481F3975D1C6ABF322F6B3069FB4F39FB07DE9DAECA5940814EE05028BCE992C095821D746980EE08069334BE9DC444C06B0AF1E0931A92BEE0688CB8C12522F5BEE6375E965B91435E8A58CD27069B8E833168EB6300904A8A57B97D6E92A0CEBA297446011CB5CC005940EC1300E2E7093411C9F620A7C9FAECC49BAC9D05F006D5187D611EB8DE265C5D7EA3F4FD96C229F50B968C903DBF08363467064ECA7E1994C99CC846C01579ED7EFBB1A972A700D020A954A2693D5A7A15312C8D92BD48E5C5367DC4D2E41F101E080E41368E11BDF6C365AE0AA2B72C4BB62C46C749584A07BF91BACB2DDAD599ACAF512F08F486D99AEA0FB17120CF7221C63F23DC5E30FB61AF4E5F91CCEFE5588222859D711816FF6922A0936CA436385D755359A054C515DBC7595A008AEBBAB3EB32F1F08E998A304D96EDEC8730F9018F701A71F278D9A0990C522DA12D481216EF7DA447CF33C8B276279EA3F6C82AB97A9FB506336A3CE7E37ADD300D17F403590D8750D9328F573C6FA43856D38A3D67651179913DF9F597D76D7FD2DCC338047CF3674D9EA4CCBBB87585C4885AE3108A0CD6853C10680E6F696CE2EF4368FB447CC1A62C04E8CE4846850A1D999F573470BC58FA18B6D24C156B89A27246C56BF0C4A1FA530DB984B6931924307BCFE5E21B905A8ED834E5D70A7A2EEDB3518BDDF02B8D131AB69382E6053754E1AB58D1503D30CD321C644F2DCAA8E41DD5B8F4FBA9B2B4864B4BE0167AB826DBDF70203FEFAC445C981821B390CED6992BEE2DFA538951F4C7BAE07CE904CD4E9BBE19C800E0F7B3A3446B602089DC714D9F316B282C98CE58CB758CB3BDBB4910085E2F7B9F9550BE643C025021085674309EAECE41E87A26C61916C45B17A669C4CC62117D1D4B9397484314012BEF35213DD6C1CE705F585A07CDD7880A676876576316196CFD757DE0F604561E38BDDB0CAB1502D9D8D03164FC05FA5ACD052F28C86F60C8B03F99E6EFB2BF79C32886F31C45644B4BED3A5A3D1498E906B6C5B13B2A4D352E276FE271981FEE09832F3E5762FF5B75D6097D158C6EBC7CE79CEA808319AE7A8EA4C199BC4D4B4FABB2578F217D8F7187F465DB85D1E7F1DE97511478FE672EDDAD7CA3CD53AED21D0C6E7B1E5C38D30CF26612D4D764EB82A39F48C90B8D009073A6E7569B80D4E99A12434072C5A5CA5D1C09D6E595270A939C6E6465D6F1EF4BE316D8C0DB45E3F72C99DECBC452C38F719CBC65B4646F22F4CC05068621B6ED1C29A9A15291696AFDEA0BE0E9D9BEBA973A0F51232FC18098AAAC28CF98AA91CE9104FB2CD9D949676BC0F112CF4336B706EA2BAEB66254572B0BA751DC9CEFD8EC59BE46F7A73F959DF1459049F2666440AB03F56A643DF922399C7F3341D0022599C89D9B9E901B670F9649F785CA1F82DEF732FCC51A2143AF0BE825259C93F239E11942880776E40110F3DDA0CBB495B41F805193C6576AE8E0ED48766BA1C2EEB0850E15AF85A085EB22C7AB42605E7C927CCE5E9B6B75361E7E176A083671928F06CBEAB5BE1C2E8F982FA03E3DD1249397647FF639E16863A71C6768A37B6AEE5A98E8C31A64FA88B5E3CC4F342D8A4F968306A41B15F38CC8E7CD14C946702160D8EF792681A21E39BF752999A93398A7218EEDD7A92FF595FE9ABF6AF846990662490D32622785C6C7EC701B4056FD87BF6263252E0CABBED4B8DAEF990181BA64E6F5F4B458C73224A3A187D3EE728A379C9EC14569D52A872AE89DE381E6B7DB11F43BCA04B7182C97BD05F4A2F2C99061DCFD5AEE67EB9C148A03AE0BE774FD8492CDEC5DCC6F9EABE9EE77F7072A031E6D1BF416B11DDD94F808017256A294B3880A4C9BFB72BF1E6A837E1B92654A7AFA24BBBC801361D82F96A4FC3DEE073F83FBEF10014359738773525E44D5287817B91E3EDDCE0818231C57ED1921F62224B4054CD8DB3CFF67E3B88C5E33ADDE2FE505DB36713054B7675E1986BDFC599D944FF85EBB0B3A7E4DB9F1FBB747A5B727180AE972EE969E28F5E26873335E17EEEA8A6AC2F73994467A05D27D45DAC549053BCFA225E00F2DC66A38629027975290873D5AFED4C4B4DCC910E11B4F3C9F5E6864C1B8BE6EA37775C93E4EAC7C0E9E402FA5A129C42410FD8E05FC33B3ABEEB5BB51EF41216B5517B107AD4B4C9FDEB7F9CF8931FB00B42522DD0EC6A9B4FF3BD8759C0264E8516C7FC30C8245A2FE67653B56D57D18E19A1786ADB8DD19EA88277D3C44297F2258806B05F742689F2DE7EFA73DBF1BA220C8DB2491FA79D89752902CE2941705F78E07581E20CB8FE4EE006BC7137428F04867EB898FFFE03FF473AB2882FCE1B18B77F5C26CC56F0E21BD6524FB73C76B25159F1E5E47DA471572A304DB00ECF9E4B87E63F8AAF0192F00F1D64420DE5A7D1E7FD92CFB1B9C2DF60BE5B0396973585A42807D4077FA46BFAC0A431136905C4FDCF7217C6EE88B4E890B0E4C2C16F8B7344983013C48CC906C1840065B2CE2E7B696D1F23CD5DD700BF3F93CA2D3303B3EA3EE5AC1455D12FBFD69DE3B9D1F84D024FACC5442BCD3AC92D3D01F372D93620B9B677986B226A945F33504348A045EEA402AF159BCAB414D72C78D46FEDC4BACB40CA2C88029859063BA420078D89AD117D4D64C59390BFD158DF792EC961A8BCC85C94FC64BA3EDBB56F4659EB475E29E6B60C8D79E69706C8513560C4F1B57088660E1B080EE20E86A92A00D530AFA67D98E07FEFAA3235E2F3F26BBEEF723F471C9EE9AB90B28043204017A5EBA7773EADD68D6CB0D57FADD92ADE229C3CE3C25E87DA7D2CB0CA3A191983EE598DCE5CFCB58902EA12BDF5EF6FB7FD2040793A5FD2E68CBC7DA044E8E070D4C00637004933A0E37B99677C9542812571AD24BE557B467185E8B08D8762931E43DAC974BFB6E7EC7A5869F407EFC390963654B8AE96E64021B19EF22ADA0B66D416715285A0BDD9A7D5263DEE4B7CCF84E39B4194ADB4CF9CA10B6552268BC8AF5B8DCD2E4C660B34884C9F2F6C047EE9D0B9FDF5E89DCAD93BFB6C6D3FD3B3F15D69FFA1F5F0638A6E76128FDF3E3B5572349C1537D5A000EEB9C8F96B31D0C33FFB2132205BAC68A1B92A887D21AD985B0B0D01AB69A4340B0C439E5023364F1841E2E458E3C390EF23FD9CA5E53AB2E53BE5F0DA3832D67428AFF8C99317D7F8E1FC2C4C2FE0A9E6535DF18518BFE905EA1DC3692509229025CDC6E6E813E99CC1B7EA970778CA59C3BF71290F5B82A527954C6DC70F959F1F68C78771313A1D70FA6F2419C19B126048DED3CFA66880C0C41EFC5B56C95F558D0DF082A0ACE6CE10E8E2A790DBBE00F53459118EF686D5844548FD83553C41013FD5833C9A919A45AED38AF91B34F5E40A8AB9F26A9AC4AEDA66352340B63009E109DA455FDC7854B20AF183D667AD3386669A46017AA3EBE1D8B19B8123D0402A7700590283B1509B71FAF17FA9AD78928F5141176503AD7823AB20D541BBB443B2C86DDD21CD97456D617F1DC3F42E5F301CC8EB37DE43F19AB0F264D0062D6FFE23280EFD4FD4FF10942F800903025129B924D50D574DE24F70255C5BB95872B722C16DB0E28D6B83BC5C9A8CE01AF9EB43A39C251F3311D84BA3430FCDB1055A4894E0D65A7EFD96A965D6E25C087C5EF9825E2F84AC1005429214ADB88548CB057DE8A513D94E538B10E1D270B2765091674DC49FEF55E0F0BF88B09015353FC10477027005705EFE34C8E83FE110D5EF65FA683B9E786A3A477CC9A0FF1FF7336BA07BB3501CD7123FD44FC1C515E0CC76E32CC937CAF8C7BDC2ABFA8DB32E7E1A7493CAA64C527B3E4AD80E418FD6A895EBCC2537FF595E2340F240A53621E2AF5C3C18A560F051029645BDF8AEFE2F185EC710108B88C97A7B245A67CEBEB24FF16A952064FA61898629DB168F6418020684B674DFF2981042526F02247E4CB47F593033D633963D7F1888F07F51C1DADB5276D355CF9234437B0C1784AECC8D8637FD9503B9DCFBDEDBF7E1E972463B4072CD8CEB5A8D4F4D52598BA33E5F57653852A1D0A070BD0A37087F71160F655F500D40446D188D118130BA20D92A13D03D9EF857BB53EB4494A8FF9B301659F1F5C959A5BB1431ACA25B7F0BB2A511D3A84515C76A7DE383D6F7D7D6608B943B0CECD8B6A9B277373BC9D5734AB2967A4D0E30C5A00FE1666ACCF89D3A341B5F5FD9F2BE3ACE55E6FF73E3056CA1D159DEFA28765B775C6D5798973F7D4346180657A7446F3836537208EB75A8E3E9A47EA0695CB164A52A9FECDEF761BCAC90E3DB02286160D350788F79544ED931AD30DC960A9682E66F08BDD0C2B865A3F2F4B8FDDBE3A901A3A04B1CF50CB3BABAE5C414B180866619960401A94D9FB420FCA61E4F5C9B647F2B78E3E289A4795B9DB4B8EBBEED4A555BFF56DB838E2C76A692CB7201F7F4C099F96E80979C7A617E17619620BAB06ABCECDDB32D0F3D474C9F208405F5F37BDBAE7E9BAC6FFC1A30E3417CA0AA05848AD5AAA96AABFB9B81037CD24A984FFC13DF3B10ABB51C53B65577F1D94CFC108941E8398E7043ACEBF908B9EB43A804C93619474370F681B0ABA24A5294AC59B1BFA00D04B6DC8B5EE628193318689EF2DFC89AA2E4E9D606D2482970F90EED889BBBF676974CF168DD95DD4037B7A64812600057E3FFE0FD8257BE384D6AC6FABE740D0FBD3A9EEF55B0D5914012CD8460A69028A0C88FA2420FD67C25C85BD1E9D64DCE9B6E7F052085B5FB6A87041D358AD87C35BC875B51D0DEB283F111F50E9E437F301608300E7B375A050E1C37CDA24FBA3823E4EDC4439AFE2DA31DB1C8AB2BC3D013A9C259E5ED0DA5173342A55C25A0825E6549609938C33EFFA925864C35B4F2D389F3134C1E53F7BEBB56869C248454E78918A879E04562D808684B488F5622563C880026C71B9285C63EC0016EDE2D1E710E894AB8159C9405B105C03C3B1D0272033E0753C7251B83E363BB136B6C528DDFFE226F9C4CCA85E8ACF9016278F52378B1AEC9165FF28E152C83D80E1481CF4A3E422A354ADE53685F3CEA089AEE3A988986CB7A9EBB153D6420EFCB04DCE8F9D26BE9A9CEA8AF8CB3BFE215A3A08F51924CB9F555D70AD105304D5CB5AFD9B173E8C55781B4D4C53892F296A86E8DB4630AB30FEA330A77C8D16A9A1A799D70D01173B2F3DE56E0D115BBE3982C000386FEB98A15A8AEC980CBE15261C56FC8E5F202E2BB6E9FBC0C08C674A8DEB5A5B4D77DB8297540AC0423B934A99615710A328A20AABE46665311AAD93AA5B996482F34EDB735E4002A17BAA9F6E6DD0114E49EC255EC29ECE707F7E25DFEFC649193B1AED90E41CA5AB1F531ED8436BD60790AC0AFE2C8D6C4556874A5869B06497993AB5EBF3C7402A31D512C9620D8F362BB79A5DDDE55FA0F415E8FF752E7A2E799C16353BD3E063B0E564A129A6B9BCC3D47CC7D47DAE13B5D224A1E23F189976CFF80EAF344FEC1F71614047B2F7A0453940A6D68AAB52206E71BC29440FBD4EE482196903AE286E3A99AAFA138EBAE177FCD6916805637F2342E84A8F1E5C487CC1322C05BD172B2D3BBFF153169D357C007468B64F7487653848897E6116264CAB80ABB23285AC1A07F4327AE8003AF8D807CB64BAD9261E511F1CDE31E32CC2CD6974EF91A908006A9AF541A756A763AA4521D029AFDF45CB5E01A6D59FC99CB40585D476CA3D83145E08F9E5389E3B7D8EF6848268898AE43685DBC0AB25F7C7E2DA0F3CDBACDC3496184A910B067EBF7D469DA6056957694BD32ACFEC87B4FD817BD746ADEEC8801F26405B911A97CF8AD2B5EA64DBC8BB89583DE0B51C4B43086AB61CC776B91AC7F41A3BFFAEBF0090F49C901EE142614F60C981E06937600724B97ED22568453093BFB9E167CCBFFBD94177F2E0D3CF868B4EFA30F4CCB1A623DB42EC94AC7519D5D2519037E34C436D991682FDA8417E114C19F439A383AE267AD733F68FA053785D9036D369A35E272747EC7BF4DA27DCDCE3700EE662B6E7FC72947CBFBF89D425F3C69589AD66A256D364D505DC6A725615902267D3B0882302196C20B77B307E449D9DD8A1118E4BAB6EBE94FD209A369A0B78B0F5A3035E4E07D2D9EFAF17A0CC6B3D7B8565CFFCED8C6590E18B071EE22C90020F826D86EA3EBB084824FD8E5B8A5CA0B62949DA634B07821AB1F4CA81A174A685F9B096650B5EAF5C1718D2F73860E746630C1C7D75FD09DF257E0FBA77613258EA955F266EA6B1AD336A83854603087DCD6CDBCD4E56C79F3E06BA52D563CBA679C6EAAF7ECAB26D3B97D265DDEA58222A0FA69F51CE33477D075C26729D58175964B13D8569CA30161AB97552D346B548D3C603B4AD9C71BECE589ADE0546E0B8301EB72A33093455BCA732EDEBA0D152E0C059DC3ABC76FC47C129C3747055C4609D65CFA5CD97BB69A15046C708C5BC906741A805B85525617B797630E95A6C57F479F8F1B087544CD7847036C7084737A1B78A86F2CC19BB51698EE91683873B9ED5C1E5E6508D063FB6C9F52257E0DD941C8E5D39598550A87501A38EA17E411027F86463C9154FCF7FAEEE4445D93B3C2E0BF312A1F88BD41263A207AD1D07C52ECE9CD5412DC47804C343EE7FBABCDDE5B66CB2FBDDB0F01490F96D620389DDE36E18CF49F196A69212CA11B333C6993321EE91A4FB3832629C78A57441BEFA336227DEF8655171C9F2BC74B455DBB1204A62A4340E7FFC546C1EC2D68441D116C442895CF78669E132D74CB84A3586EAD19EA029F2D8C17EA9CCF459748A3DD44585EE354DCD8759BCE3A0D6717C48834C52688D788268F4EB2E07F8CFE21E2631459340B67E6C72152E6CBA502547E6E0368F5D1B646A24323A67C4F617245C09AFFC709F2C5B8380368D5EC8E7A201069B8547DAFD79D3B2383343F8471BF0B583812428C29BB55ABCDD2C980777ED780CC5C22C31BC113052CE8249CAAFB6246FBB4E2759C68D89A533BABA512728C05F2CF13926056D08ABBC9229C205595349DAEA48ADE456778F3F4D8C57EE779991DC8FF1E20E97446CC24428B33AE4721673194E6502ABCC400D231465B729925E9665C7FEBCB31A70083EB8680C81EBE05955B1A46BDA81B2CED3AA6ECEAC4EEB11DAB5F0F648927703FF5216C4896DC709B6FEFB5BCFE662731CBE0B0988F87784C66077D24202CC12F2353BA63E66A52268C108D8824FCE6F210069466CF4FCF7CCCFBC5D6CEAE0E1ECB554207043D1C8A13136B64E73A0260AB7CC13B4E52E36948E47B855299CF240E0E71AD27FF1BD745814ACB12D3215FC4C39E280B6C33375316347ECDFC40D362C3B361080F827FE13FCA77005610D582C1C81D499A67F6DD670A71B52E334E34DC0525D47987847CE08B23D563CE3E4611BC1879AD77D09AF51C501D3F5CE3ACA1C1785FB443C0C49F6AE98CD3C50EB799CE24C75C2A4EF541C619D4E97F70A7D40B7A46ECC1D5C392430068038491C2D07D8C11B53915A667EC6D5926F2F889E6B21E26322A1C3F9A85020D8D14A954AB64878A34579476EF2621206C343EC2CE3E8F08E04A7123972988F2D629DA3C7FE9CEF19B6CF544D6FDE5179EEE5D17A0093F53F72D7B38EB88A799D48B2C44D0C366E8FD86E2C7D0DD7C58E8849CC3B21A961EAF77EBAD8D8D588E39395EC2C234B1A47CA91B5534A230D9656F3949D7ACB43B96BE8AAEA7C10BCFBAA4C2F62A575F5D21502E439A4A750C33788BF5F683B9D21B0531C39AEF7B450ACA9B94C9580C93533F5F4114E847BFCB5138A2210689676601CD26DF6D35B7493AD85BD61570F5142543E4BA69D58DCC64300D405A67D51683A3A9ACBB363477A2855FE1E4836AEB96C708D1C12909168ADA9A7F2815FBE59FF77E952508F49130A9DEC7C93CABB5A8E4364B1CA45E8F38CB4CC3BC70DD9BFD1BFDF036BCFC95056271B7BF7114167445D2D447B57AE482243C2951A87BBCF3FFE82964A1B932AE466BC9C7EA7B2C2A171D86BB4880BC711D7FC21227B7FB4A4089515BE46DC5D9531B5F875A488651880F0736F4787DDF8950F8E0B201E915A2C1D523AE86934C9D3A9F3F527468C64AD9F268146BD547806DDBCB00447515E645D000AD0736304C567A16983CABB182AEFE13CB55347E13CEF94C7D8F06EF39AFB8111E79DA768735A2F02B637FD896A8772FE56948211CAE105E9A64C4D06E98CA580E59371441563B1C994CCEC6392AFFFFE985A309280D35C1C3661317B85B347812497D0A595A914E711AADC778200BEE1517405194D6BD349808B508D1FA5C3FE306689E640179A5D3A945DEB397970292107B6EFE7019795BDEC201E09DD95809AA5A2D93EBEF1B397A8151769A1AAC0B39BE890F53C62B6B5263DAD4EDB9C1F638F509FE2EB8D48ED2DC9075545D6C159211B494C5176D967897C278F3E59439619875754AE0AFF29C4F7EB106355C0C437F5B74FECE36B512AC9973272B41786A536B0A481061CF81198523F39E780AFBD8CC35024863382E523EF6C9A692433439C85DC83AD6C25F84C9A50E4CE869CB76B61082F963B39A64321CDB9EC2631F4E1D206FDAB901A7ACF657BB0401F89C88442A7CEAB34DD2970553F7F942EBFAB183A703AA109943D12EDD8751F75AAAEE6F88D7D9A5B01F9C49464BE31658A8E4277E7CF7470A5E9A99E3C63EEF630F9B3BC394E09715F10D7CAB9C63750A7A0B54E50AC9CA3E7AFE98B4F59DEA31AFF55DA1FB8DF64E65DAD242ADB9CE759CE7F9E13F977538FF2CA89E46EEFDF8F5ABF5F44D9E917CF4CAFCDC610093E9F7A0EA507887F938B559C1211120BA84CCC467D9346302B3D652FE8EE07D0EB334AB7B2898C6653B4E5EFB3D5E4F88E7D2DCA4CDEA467590037E91D2D5122BF65618FF5F1BE231C9590398EBCE6BA9CD73AA6667B332E00726A024C03473CE5FF51F68118D73F825FBAB4DE38F49DC24060439E8AF56DF5EA4FBF2D75C04E448D7352835FF01AF6DDEE049195089CB38DDE81FE4B07E4C9A6F712F1D81941D1102CBB5C70F13F8AFC5B61A5303E7F56832DDB78985951E680F265118985075F72E41BB4D48812269BE2BCF90F118297127E4D6D9D1826E12EDC520468CDABBF3E6C8B569554ECACEB1923C32C20FE411F6B2EEE36782E7F0186F0A051766115CBAA1355027581B291E216BE18B64A3708EFFA91A2E70181FD2E63C4BF7A288DA9F5963FEB84A8A7ACBC0BF7518B6020C3202780148504C32B05F171AE78AF37FD4934193F4CF54B59509E98A1704E8A7AD0D67D8E0AB852245245753D0D9F8557B55491B4C300EAFB9D96846E77E53A2C9B87C8FB9542DE8D63BB1551DCFF0E59E0D83253A56D047A6FD322F2D6D0709C64A464C2D0115EA075B197C7280A6D7863F10D9440EAD9B9AE624C7B4A2612C82EBD4CA34B7DAA9D8F019E90D9BEC1F55011B9938D96C08C3B33F3C4468F76D67E5B2A0124FA3C046C00B51C70F30133AA0D6A245DED6D247B61F4039E8C0A88FB7091971FDA15C0378197D30FE546FED13996B6FFC957B19725FFF88B66E06CF8E1F0C0B1A4718995F43FEA9FFAC07E6B78D3A3266CFAB8BEBB73F351BE56FC0EFD4962C3FB890855E2BC86BCEB5AB47A16392A31CCC1166FB91251AB5893CB6DAED15EF50A6C3A543B49608293439B19F19EE9E4DDCB46CA8957BEF47FD9475D19542D445C28DC23C0C4CD6DE2B8B97866E072B9E460D52BA1A69D4161092396A24DCEA56D27E5BD0901057E8F21917257DCDE4C778AD5CE49DF7C49D5CB3ACC08571B92D0FDC8B592B4D8D7ACA8532CDA6B644071859790305A39A59C3A72A0DFD1186171EF9D3064E13A09C8B0FC482A3941BC251F8DE090E0E15C4AFE433015D45FE9188924F8B378F947F9C9677B0782D52AB6AE0277BB52C21C91536D743C245F9D6349A3F384B6F6EFB7E6517AED14FB84F8A67DC2871851CE06AA9921849781BB683444654CF65AB829CBD47EF4627407E2820110860BB1B224598620C479583ED508FEBF245AE05E5189BEF5A12383789BECBF871F371F6F6593C89613D08067375BCCD9A402658D5140F9E09A9611197363009FDFF832744B229008983A538DE37FB6F4F27F833443CCFF9D23BE364D985637544576DCBD593A5BDA04C7F2AB7E9C05727ABED52A7B80D2E1C198FADEA935ACFC0CF448AC5D99DAE17CBE3E40D9255077F238BAF4E8B2BCB160AE6826913D8185D60695F1659E1BB0DC37E73FD83D851F6571DD64B5C7D00F661CB0A4A6E94BD3A46DC8E60A933578CA5FA72960821BFB4C5086FCFF50B38BCFF9FF230A6808739747E823CEAC422C23F9682831F76C6C87B4383314BFE5FFA019BAD1FDDC86DC7C323B1D2797140B398BEFE09B5DB85748A6C3AEE8459110EBF19E7984317245B5A3C771B487FEC9A37459730F0D5CEB09E8E66DFE28B771C6AD9D803FB9A6D4C554B5541BF722814E6EAC47235D662A484101F20349533F4F0D9C5F73DBEE2C2D37FAC908365D258DEFBD9831BCF14FAB622402237E5FE81949A63461AFE455D902C25AC7E1D8FDED6D98D1C1789F0BE24134017238227176BF7BBAA6DEB14DB12E960BBD0B042F95858B3646FF5EF684AE0A6F525410DFAAAE680B434857A431359B9EF945DF34CFB28C3EA1C9859D5564DC53DB3BB3CCF0A88C01A36E32683881A556B758EFAB14B6E2394645E234B11C00A6FFF98745D48A34B0923F40C249314619FA8E31953AC2F3623179875CCB93F54DB9A2DDD00D6F0F33E8FF39B68E7A962D6BCC2577C2ACDBF705DCA4ABCD1371A0946CFBC59D69EC479278E7FF10DE4FA247640008838FAC28337991F74059C952AE9ABE8693C0B47BA447F369DDDD8D8EE76A7632396A28A6240E8EAB235CB7FEF3A5651D92C964D424DCF881AFDC4BF9DAD80AF5C5D01055A510CEAB796AB79BC653BB4B99810AD21C8E95890384C211CC5AC8CEFE7017DA0C802EE842464849D121FC89ABA6D86B43AAC5E51F7C4C078A4CD588F841B74199590E534CD349626FE23F4376FD6E81198440DD9D9DFCA6693ADE758BF0CB33D94F3BA7040BE442C94BD24FD799D8400E6D31457C8433CC1350EF3BB79EB42AFA428B9BE14A570FB58A19C1AB147A6813E7270D795EFC7798AB4BC17820B68D915B9B6476536AF071485F5DCA699053EB2CB169A4B0240C14B9165F0F1D424091374A0F07393F2D5F2E3E86561303A7AA37794960C9D2E22E811CC916946BBE925FE11F63A9D76AAEDD136DE12B43D8DA81666F1BDB5A05088404BBED8DE3172963241653824CBE7F327DB226970E4FF5156855D29EA2A09C139889F1607317AA4B4B9A4831EB213F5C0F973F244E39004F0CB0A24270F93F37B4D44BDD0C1AEE9B9B7C8E9731DEFF1BF0C64A833ACB339DCD6626A3A325047A8C1748D6BE9DCBD66D144F85A6DC9354F850B4E14AE265A61F56E37BBBB2C964E0BFF8912A4F98BE2B9E51BD37DB7354A88BCEDB72B90C5DAD7A7E6AB17D525642662A30FE8D4C980EC6D262B61B76D428E45A47AC5268AF1A44E7FEC333A001CA2A75C145C9F2F6894E2F407C2E736F5916DC788CF94A67D1AB3F04C2209580F0FA3BE349718A66426F26F87D30E606E6BC28BAF3C0D3BE2FB3CF247F70F140EE1828BBDEBF6E596175DE45A63B1D4E8E339625331DEF979AB6AE5BD29D5784A53A6925822311853145E9994B4C360359169FEBCE908A4DA377FF09DF71B3C88966A7A7F7B7CC887D2173A45EC73BBB2C5941C667FBED84A639AED6AB0EF8F09A029DC6AD9822EBC40BCCEE8D175C6D0633440395DA6858415134E13889BA94DC27CB303C0E245CA5840C53A14FD9DE4550C3FA337BDFA5BE729960025D191289065401CE4237554037B937060B1F6537C67FE815D0B20BDA52A0583056A3C36CFF38E09041C5A2AA2F6AD5E8B86065196C46438BB9C9623436FE140239940FF035DA645D52BFA0678139F03ACDC5826BE8248C00E9932D9BE5F173A65044B3050D427F49A65F5FFA09D48469AAFE3B00C2995124C2C5E16ED990D4FB651F2A29A4EA9AB196B05FA954C1C961E3D82BA3631ABE3B4E7129788A1EE961C615D710EF4E16B62B9759448F0615ED1A9CB1AF9C5BCA8BCD076282F90EFB333E7870FE9C60DCCBD02C6D9DC5C7ADA1A6FEF87C97FEA52303F658420F59A3EC4974140ABDBD1CF92863D04746648C1944085483F284471748E5CD84C88035BF9B136AE2781DFA957B8BDB018829370DBECF5D1379A7495B23F6798495937970DD9F9A527042CD82EDA2BB8011AB731C3680AA84500529DF2778D8F7E795DB4030DCB75E1A58E8DAD108CCB111C358C9D10870225E2A6F5D01EB6802CE87F2771FCF58BB615A390205BC5F36C69AB8626F7246CD958BD06790D12FAF7EF368E015B0B0EFB1EE48DB68248A46817B9945200B8F31C976B477849E24C1F862CB5419BDB6851D991F383F7E2D5DC126ADA1B55EAEFD3BB3183E632EDCEE82766247E2CA8AC63129C36C8C06B19F53940E5CE5C06288A1F097F25DC52F917002145117F2F791EA21E9C3761C314C59FCCF48F7B580450281D878BCA0682984400E207D7284537A56BDCC71B6DB74C5361E3A521F38F031956B73C9C11208CAF0CEACFF4483AF6220AA1CC822EF8D44F219E41C8F94B711C5D42843378AD4F87294AB16A9A88C29B7DC3FA8A8E3E5147CB6FD1E7311CC42C225558E5576CD4FEF4D742552C535658A1B838357985B11C7A2AF55A8D18EB42C9AF276B2E264DA1D439308CCEFA183BDA12B78B9A6D59C27A235A92E4D227091E5BD43C9865768A4288C1C6329BA031F033C96E91535B2D82A691C883C8E0FCC7227169C50E18A413CC69C633E488FE7DD16F7954CECC3B724DF579A77E88D9B41C1A69DF51FA3C2F75B8E02A524D88A135486ABCAFC682D800B9AE8731EFF3713D92EB7C870393D23C7F3C5C49A13B039502387ACE9347A96B76E11DE3A198B2B08EFA63A8FE94941AF8A7E6B112B194B853D9C9008CAEE337449CEDF3480F791016C5C56C71AE2922F88C0F96684A7FE2145AA2E3DBF70689ED1D12BB01E122924A4A0EC548664C5EF6B0B646493AA22B9996E0C1E4FB8539ED60B418048281D7BD03C642C18BD50DB3B9E9C3367C4A9787224D79673889698A02EBA93AD1B9CEF1358B3990A2CA17F166A5154D2A1E24FA24774E2B08F4E414E7F01B134058D631A54A444A0C6CB4954E985BBE5F7FCEE09BCE5C8410307C051FE3A3B1BB22684387F60131988AC5292BE1547E623D0924F7B01893133E1BB985AC4AA7F1CA6ECF2AA2266E7CC22AC3BC2271755F754267533D448D3EF7D5913E1B8D63446CE1B28B0FB19705C1CAEC630762891D97B323D2215E1A13E5327D5A4BE114A3051C4BE9B5BF04AEF0F95914BBCBE851E66DB54EB7BA8A1C980D0F2B598BB93D9F0CA2EEB65895191E8285AF6A3ED832897495A227E73A57A56ADF1D71A5ED68F06B962AEA334A873A7EE4D54A4A4DCF55857822C3652E00F3995E4D365547158B6BFC63607A51C2AB115C6C7AF5734C5372EB404AEE61DB0653743181752B03B15739F23D9850880B5C82F59DE4E26A01E46D2DE5AAD2A5A01151D96922E67266E994B726DA127A037118C6E165E5240AB3EF5F213E5EFDD79D07996C645E6910AB6B7E182E2751D4EEEB921AF71A1A0738A1CB2DDA3E4938C65E109AE4E0E8926D1CC90998F54BCBFCC596B6CE024C262C9FFA6EAE2A98FD831C0558B44664374E768E8B6F31EDC1B06E2B17D7B981E328F352F8AD81F08E731F74B19805BF2B8DB3985A725DBA6F140C17207FFBA28DBFBEA2CCC34FEEE65660D1664CBF730D2FE655F78F79FC7D707FCD1FC2A5BE199C8056BE309E5D3D0C67D82E1EC935C70B73906B327FCD7B403BEB727721ACD9029F22E312B6E1A24031725B521F29E76D75EF1043F8992496831D6B77E5516160F931853E49D7128BC35337DF55FC6805F766EA9CA73D927953A353AA27DE88D0742D529BCBD431867EE09052233BAC20BBA48912F13EE8AF2A0EA9E294CE6EB0AB9C3E3473366B16C72CFEB422FBA8716C3BFBDFE688C50A7EEA8A4DFB1EE6FFA37D0D3EFCFFEF507402FDF74D3B43B0BFF06C5E439959C0B830C334AE9CF8D0D20DC4B11DAECC6F0F79F203EB56175C8574995DD55F628FCBF6FE8D11CB1DA7E20D7ADE37EA8E3B0742EFAE94E0A08A95C0CEAC1945965914FADF7E973B1102B5A6BD9810536761D1A3135BFA73B81A4A14F8035DF0983E971FCCD46587C090D91122E313E46007E7FDF45BDCF808B549A77124C330C7271CF74142AFE27CFE9C75CC37815BCEE5ABA087E2F939D4F3CE5E557ACF21EEA76A1882AFCD523D76DCC5E9AED83D07000171E7F971D9E29766956BF51603E660DBAC5E64F836BEB89AE53492D26E1B88C1F1C16C07007B4E731BB2BE3C5B4A1C09A31A4A50B2EF34D514F267C251A085BD5B9CBEBC5F7EB7B3E578196E4F1B4E2E50B8AE2A11CA7807C02F874E4F99DCF182E8FF94A05F9C22159E2188F24CBCC535CF21E98B7CECA9F506242F10A024D6E9E03CA9C58EF249DC92430FD25F48918540B8C7050EB0A899ACD6F6AD2E04A8F381690E595CB4370CDBC5003F1BD04500FD14B4D64291AB4C7C8CE70CA3B942E66CCF7BD609717FE07F1974713C75C4C9816057503D1A49C629C55A540F537CD60ED35CE0F0D9998A607DF9E32FFD847278BF61EDC4061D81FB38BC2E2EB1A41723252D67D25C73BBED8AC0DF3C690EEF5AC9FF651E4006388EB6035F6CA368AFC928599E68F2E89AC830B878810C68ECF6AB892ED99EA093CD08A1F7E1035F193FCFA749997E3D283B594223E9069B5EC45F561FDC9E6C3EC14B65BC5F1570669D611BE684F04ECA0473AA8DF8604E23A6541FAC19731F3395E79D5B4C7A93D7B8164CF3BB5E2CA8CD0C865D0826C700B7D35B8CB250608040B26FA8D04683038D0D262458F4B70F855FECFD1AE223F13BBF8432BC5CD8015060CD63744E1EC1B454748426BC12903229140F9F8E798805FB34A6A9FA58566D5DF2BD086866DD760C2D92A344EBD4C2532A57980D4117766021A6E0415817023E6253C96F614A673BF524DA60B63ADD0538BBB369262995F5FEADF8AF592A550EC8B5FA18354868CF858F384FA25AD5792FE0C565B22F977A07AAB000C48232165435592CDD10B481CCDBB13344220E665A4B30CD35227EA736D049A04454FB459C79695762FECC69B7340A5D0AFA49CE0B69FD3E6F2B746C3678BBA12EE91B7CB4A16BAEF5C99110CA68A159264C2B31D010252094EF52F008AB6B250E7711EEA1C15A4599EAC63D9C5CE209E881D54A7B78DF3A004698DD7C45F91D29E1BCEACD919D09824DF281B3F5E9CBEE1D335FC686D2555404CEAEC0C6CF8AF1170F5139764CF9AC8F1D45A0924D7309C32AA51C4E015A5D0A52F12C919B4609255F36C592D483618F1F780FFF4B6FA7A4AD96C71D7435742856AF450AE241CA8C7690A8E770E893EF6F2CC837E59263A903E99A5E0679E8E79FC385479224EC8935EEBD32B4F1F203218E254BB638915ADD83E5D6530D64B7E3BE1350F30D102CE8A5EEE7B3BA8026F9244CAA7A13B2AA93B4110E79D7CC0B1911C278A0EE950372FE38B7B171A9FEAC259C12C56F20CE77CC02D321DA89A2EE5FD6344E6DDE08F7DE25309C38CF5FC96671C6CFF116864CF4F22CC1C215DE2165B1B2571D90FE8A02CA5129E517CEEDB2B725AFC48DCAED2C7179D83E3348BA6B8D48F50A86086C3DD7967AEF92BFC502C1C95C4AD41E8D74901F6EE0BF9A18D2DC284F07ACD92E6414228E381C31D4DEC8DA2D6AF6F69C8630A1A80242BE245F14055C85D8F81A73628CD6A068601826193E438646F622BEC268BE9FAA8669C9C646A2CE46E25D20036B1A9B6EE8FA54D4F3EE9662EEBB3823A8085312538479458842C6F10B89282CB885B45DAE48CC7D29C125A80ECF5EF370C7D3517E3CB986D8AD1957B29DF9E3DA16536132CB52A10A37C75EC945F5F06683C49EFE91F60CBF9261788CD13303634903AFFFA91964242C808E6DBF06257B05ACF87D5FD534E37F77C9BD3593085DF9C10C927E7F9BC65C7292054E871403F36FD973BC24099F7EBA9DA3FFFBDDBD7F409E89D3D745143E1B6E0D2D86204E76AB6E74045FD44F69727130B841AD5CB9C57921658B5F7DAAEE29B346CD324918107B2A541DA93D765CD388200A679C908080093587328B97EFCB79B3806DF8E3F15108EA771E774034D03D2C99CF6377AA65C4676D0B06BF56CD433321A522051DC4FDFF695BA0615E31AAB97CE6668D3D4491BD1AC0251D762BFC8BB141C49F9997207A0485C4C2E41F59C7B086B88AA424E920B362FA722FF4DFE8A0A884FF557936B57AA64527C8F227F19D895D3E92BBD9795BBD477025B592A357F04459718B19608595D0D4BF2D91F2300CD9A279A3E5EAFB9E4E7046ED18E5B4901A65C991563CA84B6B2FA6A0F40084B1E941DCF62A106F88011FED5F2B2F1E0793E45B41F4BE86DF17B71E1A8E5BCA147EEB45AC753203911C10CD36FB385718C66952091B112D19A0CFB5123CC5CF55A0550CC8E4D6AC0985701582A0D3F8E50F20202A5620DEC7D6E49369B44EE1207DBD8D9C39F21AB244441296D6C405E9881813BA70B5D5C360455C9A49EAAF65B40669723EBEBCCC61D2F4A645D86CADE83A1CC803A39921C582F399BA9BC6546B02BF4888E5383F4086687AC1C137814FEA07E888C45FE014CD2B1CAF6CDACED9B0AACDE21FFF783F38C2D1EC3A183E95B1A409A01B4008A626081026BD8D2C830D2BD5967FD53657030766EA1F47E36B7F49DA79A236E301FF8F4BAF5EF123D6E28AA69C3CE613ED93CFDF8C9BD6D2AB14C12977AE038AB22C1AC55CE2A7A2FA1F15F0BF61885949661FF05CF0FA93D3949C9C218A26F72C067225E5FB66C3568269B027457BDB78C2661118118F80828337930ADEDA27ECA832297FC47E93A7A2F82BDF71C930D689AD64C1499110AA240ED1E09750A5EF86B44546888A300D9D2C09B62C7F74FCAFA1BBB7217AB2B62B3C77EC67C0277C247472477E0222E5B443395F6F40587414AC761FBBA6D9602197C684EC2DF2E755A39F9D6F5F1FF980101F8EE5CC9B41ACCF70CBCD96B319B7ED19967B02EA5BEB7345349BA870195790CB9AFFCD719FF76A008854C6AC3A59E651B06DE513661C186288E2B95B1A8F621EF33468C2F644309E01A4E8287B575947514F7F6015027D823D163DE7B880379BAFE68137070EB1D2F37E1C24B4704560D7AD8301C043F1A32912CB064953E9FFB88BCE34D8894D3A0AFDE4CA88A5A7B6D3525BE71A9A056BD9F1F5FA2C79D141A2B547D9A0C6C3CEC1140C87F2F952CBD1A5C8C98F3235F86F10B4C9F80D3B66422BA9191020339341E44258098297E3B7171FE9351A8C97C7EBE264FD9E38F5A2AF3A592BA48E7D63578173269441EEE97428E94A227FCEFD43D09EDEB2255237CD99B674244144A9A6610A8C58F408424F8DF0E9B7073C4535A247AA27B8E2CAABEA04E1C76A0AA5838602BAC2443B6817EF26BDD608C48416034723DE25F6D7AD43DB0464FC4B0402966FC46B70731A624C85E09C4D9BD585541E57C12FF405D405040E5F702286FF56A11F0872D72B22A7836E45B657A72C6254C655B677301128076557A8BE2CC83BEE96C71A15528FBBBDA6C343FA4AE841C35228BA3A475C50148C8CCA5ABC922A03D3B1D7F91E5997FF07C08908B1C2E68C90745129049AADDA531930E18DBC05B4A69D795198880F37433DBE3461C3F809B8E134064CBFDE5062ED76BC888850D4A60C1BD49FB94119B75E6E6AAB83CE1219F3AD8B7DB02F09BFCBA0AA0F40EC3B57C02AEC5F77C0B80578026DBA19F31262582D68CFA5BEB431E83AB9DF5742A27F42A27640F197F778C0CF0F05368F90E80E85D9864648BD96BC67BADF2E2E818641D39234B84209CC040AFF2B2F17ACBAD8D0EC6B20042011878982E4F192B2B1C8762CDC19DD513DE76C9BFD1B049DEF820E599E718274F0A876DC8A7BA72DCF1F4BB07FFD31C54AA47D117C1192EBC7899AC8A6D2BA097DED71D5C6CA4B1B5F476A970038F8CE61E411B7F30E8C0901504DAEA8528BF832CCB240E4856DE317C26BC0DE643167780B79854C7B3304C3A097185F95B3DA30AB75BFF065E525243BE04BB6D0327D506FCDA9A8D422A08585BD4B38AABAAC795F7358F700267C6159D8A7CF13080D70220DDE52A76FE7965D38E4CB83232C8D4C03E60A4F037552C99B2437BC8A6DE633D84310356DEB8B8ED0876E2110C0D1855E573A57A4AFD9B0EE5247124FF4281AA5711C25923397F0C71EDE683DA3C738BC8A1EBD12D93A614A56253C7E989EB8EA36E10242B604B93009E353380720F56CA402A2A2C5B540804F4662C18E9C1034B6855FA786D479CE19506B201B2EECEE0ED16F0A1E46257D1D8FD302B80B8EFABEA9F2A1D9B8834D99CE65BBEA807F7C3523A654EFA22A319E0219EB2EE4C3F0A6E960B7D7F6EE7C6A77F6A5F6A2F6756C0A3C1B1934748310CBCBF385F4B2D268C07EE2D77F541E3BFA3069C96582AB1B750BDAA70D80860B4BEA8EED028E6E90C4D57F4C85D0D49AD53477D3147DFE9832F7B41D8DB67A9C77A481541786D56476E5B832FA6F9F2836B37CBB41CA3CF7CEC60553F3B22D4467C6426BADFEFA2B5020EF8AF2860E4E7735748C7FF8DC77BF7F8F4BB423595047145E4033F58B130E929E6FD2ACD175E18B2951FC6461B0244AEBD8FE53B25529BE34CAB5AC831ACC12D2937BCC2A4213AE3DE073F82A49BFA87511D66C936CAE1E45E6FC290A53C03BBA67DBED99A428ECA7230A40532FF49C1E38AEC6E549AA4686E12427707CCF321AB5F1FBE3FD49C7CBFDFB38745B76978218058B2E54C3F58F18532B5EE08DD7148EAD67DD04BC976037A8F0DB430DC1A715EF1C7AC25ED142101691E49F156B7C663DBBB0D27DF90434FAB660E12ACC9B3F1CFA2C1E785F486403392AE083E2F26F3E1E514AB73EC0FA4BCC1CB8DFA4243EBE665059119B523AD8D9856BEA3A50A93DAE5633D4DDB8E08E4D49B333B3C5696396F74C80D925F47635EC8C265E2D57420B2F6BB5DECE8B775CC484B0FABA661908BA2283329FC3509D40B9F952C83DDF1C8399C7A04AE9570D1314F70911818A76F9427F2BA39136080C7E17CE13811160B5AF31E8F6FA5B7D112F46EEE7EC0C14555E0E37ED6A8A370F3BFB44D7E6F8F0B59B8A7F00DCD9009DF7D1E1B08C18B2C5E003F2865FF63C2CA2F4E04915B3A09F9A9540C1D9D066D2DE6EE6A1A9DF494ECB01F4628AE83CD5BD259AA377F38DBA56EB9E60DBDAA6D1BB150888E31A6E625C069A5AD7DC0BF35E189BDBB70B2A8CF51282E6761BDF2890C4F58E0FDD6B0FE825E19A74DF1FA041EEE0E40866112D0CF18BDE8FEF6D37E0539CA7C414C285B17772752B2145FAD5715620F48622607DAE6CB55736F390B9E30984F410D89A269A7BAA8F8547467732F7B51FD496B71A3C75E234B7783592BF9B7A514CE0BD255FFD50F7BF52EC696FE0F9D73EC77EBB2F222AE8FB5CF2E9D3D6DF962A17476EEB7AC8FB3FE4BFD295E06B9DA225B3710767A15DE7CC22B510EBA0B1F4984AF7A29FB4EF320CD3D00CEC38C63C899D7CACBC059C89C9F861787733125A1C6D3514921A61B942070EA454DD50F85F0C8D98DB2C1EE41F97908ED2D6C8CA6C7873CC2D0E254AB146A158A26963D2B3F149E7A0EF07EDA5905467508507D6DF1C08C9B1064DE682C0E5175E39A2A144B16688F750FE3545853C4A1F9A803906B5FA6C8B79916E481D2CE857B5FFE2D5BE2C96C8E6D74FD8B253AC9C095A63978C2E4D9B1DA7B55DABCAB11ACCE0EC5A688AF317B3081A6DB164714A442622478EF057017FA4E9496795FF978FB0A4748B144D7DCB1CC3620E4A7D2F0F72898955F1485196A3E0B104CEC00037FFC21154E6EDE5B85BDA1D2069FDF31A81B4060A8CCF1334542566E4EB09C868AC91D6D1E7EC206E60CF3C25F34DC1B0D0A80FC69D8320218C5B6EA9E329CB3A7CD35F1C45891BE567C9FCD3A1E9E171E936B28E884DA7AD15B948AF10F999AC1FE8939774F05F2883074DEACC643C335E46AAC01938823E9E4F20EFA706FCE2CA3AC643B46C753B335A40C86EBF1301473C7BBB6D86DD9B818E3D743D54F8774F75899D2B549DACC303CAF49AB85A46C7A255346818B3CFB964DAB323395A412CF9E8C6A68D8C886D821FD3B943DFEC448C4B6E85ACE9F523117DBEA8E1556346FC26099110EC15CE9F51422248C14375EE9DE6C1CC28FD37F55569723476B2B4F253995200CC2D8193A9A0EBDA262AB239175755F42619110610A06C7775BD8413F09D3CD5667889A2BFA95A420DE341F81FC09704BA004630E2C46446BD408A67C6FC447908AD021B269693D322644A4CA0C432D59FFCB291DF48BF387B442F9363C4A647FAD8BD8335438071B5B6CC2322270E2FC90A14CE991DA6B9CDC589C0B128B1E87FE1010967FDE506457C4EBFFC76B6311A235628E1DF30E0B019B06461A7FC0DB9020097C4A5832D73BA3CD0B6DB8FD4F2E240D702CD9AA56600EE5987D6C96CCE167F9D0D97864B995B18B098FD3A6D52B496BB46B7FE9653CAC8096B1287E0E335F9395910D35DD4F2754F54334D34A26F0E2F7552E8559894E8A8F7823A057820B4D461FC04C0B82E43B7228B00966A6775CDA1A7238179DC197646AE87CF3B9E656280C82DCC7CB63792B1C77ACFC697D9E35E7ED9E07CF0BEE06E7033C549D1DACC0B16AE2CEC0F19702850D333ACCE39D24AD11F278D27286BE5EBB6A9DF53DB9C36470AA64FD646FEB35520ED542D2290BFAC78D694B1637734EC4E0A30D1351BB9691D8158BF41C151D619D13C98469EA9D69B9FDC7034E9B7D2B57B71770BB96938B4ABD976D4FD7C5B46251F2C2C3E38284AFDDB78BF2461BC4668F3F43C3CAFC79D324FE95A41F81A052DB6D452E2287F9A7649FE62162F1310A1A7020425657A028522BF9B042D3DD922A57C2E9CE730086CDAA88ED1EE68BB0515015E5ABDC6E4F30056F5F88B2BDCA16A74616C72E81C3254A1203DF025BE340DE5B0EFDCA10586F25FBCED0B6D7905FE480F0594A68628788C54FAA44922B5B40EA94E6FC5F6DF6E0132905DD4A454A7011C8CE8691560F1223C79E1ACF91DFC3A62470E48112D13046FACD0FDA80A6470E36E207736649DDABECF1F4F7E44BD37C3508C5BCC9F9E775C14411228002AEE81015C1167EF3C4C5A8D397712A77FE8584A0DC85CC4BC2F33D3BD292279617E77C7A7D3E41FC91E625D394B0EFFBCDEE0C9FB13F9DF3440F43323CC71E46E7ACBB8685ED0D9B775EB04DA13321B8AD4518B5E2B130CA15A2B10712D385C16FFE287FA43784FD7F5B5819C8AC220775F284426D016C6D2C41E61B6234F34F342DC835D4FC13D01383D8C25B49A4E461C0BCC8B212077EF5056816337ED029B9FD864056B214E9C4E14CDA7F2ACBBEB3FD136EB67D01C8F475313346B074464B177BE93006C0F0C9602E7549DD744A9732079815844537F885F388AFF33B1A86858637F40842499E32F0947011CB65064E235AB2C897ADA159AE513CFE4914B01EFD0F6D8C50E5B5863B8E5C606AA6322F023C5F07ED0702CC585B796DAFC9014B55E5207AD95928F581CE9225286043ACA4AF73AAACEBEED9D58C6B12006D22F7D74AD185243125DB518BBF887C9793FC9E0D2D94E3FCA5737A28DB75D63D5410BC1E39400F4A2B79589763F9B8AEC0065AB7F268EC9AF9B30D1501925F067A6F1BDB53C904B7CA94B04941704A8508650A530DAE2D75E9A0D330B9AC51971DF121D3037B7AD0D944972FD0CA0F5D1702F4C6B3691147FDC82EBAEF2CE2CEF296C41F861C80C47181D39C4A726595162654473AE0C8D79898B1755DF7AE0263316B1A62D085173C5EDDBA1B151DF741E0D25556D5590E0E69D92F4E8AE8F850156ABEBC31832B28A5383EA9C01BABE3485883E5A0DDCF4B11D65A33B10F9DC40A18BACB7F1059C9E38E87B0D8866F33C9B05EDAFAE956B90F0CF1E9CC32904B44FB50CFACA03C6769F946A6EDA79F6045735A4E1A0D7990DC03D12A740AFBB692EFBB6E11CAEC28F74E689D94651072563A797B676EFF5630E340387D7907334B30580FCA97B5F71D32088484AC6ACC6D22F8128E10E84B26B03789A61BAF2DFF9820C94DFD77C6BC36DDA87545FD6E4C21B77A4B048C81C6BA88D6EE95FCAB80177353C733845F0D80E129CA3DD970402E0A21E6C49C9370F1882307DEDC7A94104FE1516E50FD20F0921C199CBCE9E7BBCFD0094959B84AFC2C8616F420A1FCCE06D4A572979EF3374E85304793E5FE9B8A1A60E8621EEB099CA041590947ADDD70C17425358242770C76A591DED2F794C3B6C49324858052D45BBB60DDD5C707D048A2C91EED40156F5F718F3890033E45A075FCDDF66098A167B2EA084F0AB490609625A3A1742012D271D7C785554B05F161E6F25008D07EC5DA750C6AE2CBB14449CF78A3736A4457D786E091622D7452FAE47222827FDAA7BFD5CA3C3AB8CAFB6495BE452F1A31697EB4E8D7741C368AA0BF3CFD44BDA894CA9CA3D71A24806D07FA2862A35F4FC298F521A467E7F72C598E0FCD4ADCE5C313BDA2412C4DD4097A54531777DBE6A89E9034FB589EE4CF7418A88EF73DEC4D529ECA07FB47B5712FB7CFCDC4CDFA611E2B653B5B1ED27F0109A91C82E5107123C71368EFF966D53652E2D8981B2550AA085451F51E322D46D1722F18E0E2422A440BE95C7D689976F880A98820096B9E6AC7E5542AF473F46B6A4C4EF77EC49ABA5C5E53C21BE598B11774B94EF8202687ECC98538F931A8E99630F541BEAAEB470886A0CAD6AF69A7D6233514D3ED219C711A7DD49C3520308311FDD3E81F9EF212827ED8F55FD5459675926CB73D183373004B061033D086DA0C60914FB08BA130E51268805F0FF13A45D8A950101DB549D3B8BB81A0942672A79FAD302661E0C24E86A932872A0CE388DCE72FE89C7656CCFBAD330D9EFB0175D555284253CFBE71CEE176DE373B0415035E1CDB1D1B07E0454EC40E0A6EFB9D061EB46A8CC08774033A474E44E982426CFF44E8A21DB4107248E76504EF625D42F4260A36C15E77FF3B7C8CFDFA388564A741E5F4E47FB47A64E8F13BD29C999783E3F77760922FBD876E69C5687BD353E834A4E359EF0D7BA2D573AD06699136D57CE24E5194EB72D8939B6FF696E59AA1E86B56D7441FD9864F551CBC18CD71E010614E7CA504E55ADB28566AFCE0011FA2C8FFC4725990A3A1F2D653F936324B2F7BB5DBB674C1AB696B0E81BF0CA2FBF9AD04DB38AFA0CC4BC5FBCC87230AF6217BC21371BB6735DA5817B09CAABDA8A634573B1BE9C92D77015BF43E1ADABE9'
			},
		]
	},
	SiggenGroupItem{
		tgid:               2
		testtype:           'AFT'
		parameterset:       'SLH-DSA-SHA2-128f'
		deterministic:      true
		signatureinterface: 'external'
		prehash:            'prehash'
		tests:              [
			SiggenCaseItem{
				tcid:      8
				deferred:  false
				sk:        'A1D2B4A832DBF4A67A2A9410CB524A0596D8C25F647AFDD8D38B60F6E8C5EC00C0CC2055D219E7FBE3FD21D24CA2D4588F2D82AAC501FDCCE0B7EF9E9730ED96'
				pk:        'C0CC2055D219E7FBE3FD21D24CA2D4588F2D82AAC501FDCCE0B7EF9E9730ED96'
				message:   '296B9781103FFA753AEFFB8C42ACB3D9F5DD6EAEB7E9DF9AE3DF868D472713AC43F7AC72BA4CF5B802510BAACAD891692E043DFADC3982D6DE51CD05F7FDC7459AC565D316E2DD33D74BE739BFBDEBB0E47E8B0F6DAD72A8CBC254987FCD03E98BCA68B68976E7B913AAA84EE14D9932E94DD2FAE75310027BEF49FE9CF0DE8099C98758F0D5FEB77872627DB0ED9814C0F0895D4D9CB21223598B882D602B7528583C7A62592372AB1F979966335B0678775EC76606D9D543E9B21447A9D7100CC8B10CF4108B1FB8EF642672F6FCD56ED2320471373DDA65318BEE79DC620F460A906209C9D9AA7BD0FFA4E13E06CFD82BF1A9B91D1A9C2ABBD6CEBB07EFB894456579C5D4015F7CEB228CD468953BFF46F66994F655AC8356370B2856959E5CD40D777A0615CE9585A00FCA9EF262C7FF2551A64C8CA1BDDF80DBA297E41CFAED2AC7CA5D3A24979CB52198128C0431DAA20D73908B879BD8D4B42BAD6A4BA7382156A2243C690D98E131D328799194AB890DE28C551C43CDEC07C647BD79CE894912A320B0BBE7849AC8ADCF5487DF9BFCE82738D4F04AC57752E023EEA7608F0028AF592C9194B046B67CA0E2BB1FCC2BB5EF1E09CEB1F96BD0B2446B2D3B1668908A74540A50EB06300786EAB69629974C512ABEC91F8A9C03637D7D9BE14D3D665679E4B7187DE0ADE729594EFDCF4E2FE04D7B787DBF096E2B6C873199EE5961D4E785E4587799CDA33C8829F9C870EBAE16893AAF114EDC5D3D2FB14A83E9705253166DBBFC456A882B8ACC9B66AC5B1ED2B4825EACB5EA5540E19EE221F82E082490A6238EBD6398E8E664FCA31D3EDC11D343B1F194E2F939FC7960DE536F8F876FB8A5886CF1166674F38EAF2451B9417D359088B577DD352F9080D4CA0DDC751321F5D780594763CB6769711729CA7D4D2AEB30E4A2A8648F25E2B455E2CEDD65A6D8EFCF076B6965742B5EDC6C5B1144D5B698EA421BEB11C4DEEBC3ADD8F7C545DE733B0F5303C2D672FF8EB9296E11A6612DD99422441913FE220A2E40D774B91805DB6CB8A6038F2C0D8635FE0FE7E81903854DB0DE4AB9E0F3B65793EEE3F8358CC910562BA9E67A89726DFEF906B4799D1C23D0A946E2153298618D7E199E7A852E04C46186362756F7F6C060EC785543D5AC8D5E7E64918E71DD62D13C728033CEEA715BF84F49AA824E0DD771870FFA33CAF099D2486FA060BDB0D0E1A9A504CE32E8FB72880DC64660A7ED04F24C22AD437AE1764E65B6E5E4E30515900A293C12C9BDA9BD3EADAB67E838FF558544C3C660ECD3E11798EF92B8B036B92E2E98A6428A360FE80E304EC38EE755489E951ABF44BEA3D07F9D00CC92CB6EFC6FF6CF8E47F31B5E820A1F8FA360B498BC24831F322824FE26EE36A59491F32DBFF124437F126D21B44CE768BDC9BEB642945E85F82DEE933A4FA1B415CFAA6973DD596116F72C1AAA7B4C20BB5E4EC7A24C753FFA660A18533B3BAC2D179D016DA3C70C916102B8D359EC034641CE75FBCECCB3D1180D3BE9EAC219AF0073977F92628AD44A966F00465708A2F4031654EBACA1AF1C94CF2D9C5628D002FE2A618FF749582260A8707CD065E73AD73F12931CAE2BD52676DCBAAD35F206EBD0AC3E42793316AA7099D876D6937089DAD1492EBCD3AB69A3082A5F0293FA80E65263D67115A8884150EF5994792FA13BBC402F73ED3D3483AF5821BC58FA60F36CEF0534AC461B00BC1CFA082E19FC2AE7B7FCF4EEEDD6579783B731A9455E4AF888AE755988F3B9351D60C495CC066789CA02B644597C1B655EBCA000501E1DE08FD4348186F5E96D414D6A083BB65423B881C7623ED9CCBC2FFB4E7261FB828869FF4B21291F0B9264F41E26384B61AD2F01FBD3A686E0DAF55DA192884E626073A3539C648424B3556EE91FB4C21AD08DD6C1C45CF52BBD9CAFA54DD360014D14D3E8531BEF84F1C557C9D2447C8A9BAB74F2899C76345CF66F8BE875EA0B1E402D9B3F5DC54580605E3B9052212D28981B38DE7F417BB0134618616FE44F01E71BF471A523B6E35371CB172647A20FD0FBCDC5EBF339349E416214A998F22B7662D7F431FD2466E024D2B87619F1755AC2F96210C563BF0F256FC9899607252A413118BCFDD1CA5EDD8A4FB2495A0D0BEBAAB1BE1D6DA77A94F203C882446A738401D127FC610573B77F7D6DDE530228374CCD007BAA2B1258151E024582DE5BF72D064B834557B9AB2C684880008FB2F5484B619F62A18A4C546C541AB0A020C8FD6D6E05F77183AE6C631D347867C56938B2E5A2A659659C0C42F4C806250E4A9DC1E7C6F9EAA72EEE08F8C83D968F48355A40BEEABD89E53467F09F9F71B6652B5ACB08AFFAC47871D060303E9903FCE29339BC8A39A569C996C0BD6318FE4E383661419371DB6E16CBF78F26527BF42554B89DC0EF9B8D9C5F798B69DA43685F8782B98E28519A31F9AB26C641C842212A98A7815ED5BBF0F06AE50C0D68C2F1BED1EF959D1FBDFB3AFB96AA8C7D06448698D29D352730761857AEE64DD42D9056B344480DC8B9FC36DCA98F4CD4489E5032E03AF819A50319FD5E571CF3D8E38AE27ED41C577666D2CBB6DA2A4A7376AECAD925B8B872D587619F842F8CC8ECB7D4D9C04AF6682A5898F26BEE2C64B9818EE3E4E090B764A3C9CB8581CEFFC537A5078E03F50592AEB9B66F1C159F53E621532F51FF92BF62DCB54F8917E30E080F818E804ADAD4BD35E3724F1A415819559D65DD08D4B83387D9DECAC2C8922C058A5D6EB9A88386303826B8C6463BBB7F1252A91013936DF04728CE6105F55C9C389656FCD82CA74676F19C41A97AB0A73FCFB8242E659BE05A46E550CAFC21D4686141F7E3FA4FCB77D875AF74C7362D79995E27CAC4FD798D3AF727F71E1EEBA01009DFA829409EF682E92BDF291A516DDD6FE9E8C2E47241E9202499454E600354D88E19A40AE88247E9AE363E62AE5E906D467F2240799F2384B211C3E5E031206A41D779E2DB24EE0C293C8395C69B32E87E267F816E96B008FC7F2ED68E702631CC04FEE0470E94C60090D72AA71F04E1E852550763EC6F40B8C1F16FEAEF9D00662BB4CA7D1A3BD32EE36DDDD768CAEDEE19C62C718D5D80CF7CFB82E2C2A96E6EAE92710DF3FAAE7EC694C06D3FBDB343D431945E0BAFF99DC1BD78C9B99AC2A4DB1C941C0DC120AD24372086FA428DF5C53C7C854E498B43AF7FCF13A8D3B6E71BBBB0CCB2797F51B6E2A897F3A81C91D1219D7081DD5F8BE947958D13D690CDCF142F17D35F1662ACFE62ADD5748B440DE2EA38A086FB4AD2842BC8DB2C4F19907D0C7EED2A73BC593EF67D28310F140F71BA62F0204BDB931C41471B6FA1A27B8ADFE5899BB5C744DB58EB618E6713CB46387CCECBA46F62951AA3F2B897B22A580B8F45DB5B48EE882E948FAD71ADC033FFB322CBFA871924C0E5E3A450736FE799D33C2747CAFA5A48C953BE93237BFD47422B0799C42C48B68DA555A23652815222D1ECAB07762ABABB8F26CFD0B1663A86DAA3F4C20A6AC0E72EBEF5B416D7F0228E4589B68421E61FC9A42FEC2FE44B9B0AB90D43A3E0675AA32F295C4A8360BE13FFB4FD014540E7E698A271C56316571B3F387695042143428AFBC409CCB76C16F450463C66DB4230A348C523A9E49EF4322902F076B26445F163DC88708B2E5DC61BAA020A8A444128ED48696734A667833495FB1533329E5351C7AB1C6B1DECB12D584F4B2228C7241823A851B796B80FF9F38D77E08B1F6BF524335269594B959A21FEEDB56076C10CDBA0529D947784191576B6B286D22B4505AC98EAD400B87646E52F1BD22470AA3FFEB2B66571A2BD1D276A12C2DB805019BFDAD021010B8E57B80F3634A2407F89788E06234405E07DBAEBE08E0F2E551C64BD13A4FA23CE05D6FA6B511F770907F822F0319CB4D7D27FCA44CF106451236056ACAB4878AC69BFA3D81BD85F47FEBBF1F36152B57210695B1DA68C8DA8AE1643B06775C4F9EC8442E60FC5402E9C71D15DB913686610BD2170416530ACA6B29D5C06FCB9CF18AB07C9B8C63032D99C82D739335B4C7349AC2045DDA4F34EFBAD3FF71ACB1F480A901560DBB0BDDD674DE5587EA853F29577D11B01DAA9C067A569840E992782DB56E1874DE2EA1BC7221F86645AF365314D91414DFA9EEB186242C5CC850087D349B3720D853F27B91F15A0C5C122A96A35090E20FBCC8EC8EE0C8D09A33ADDC3E54887045E9B3B5CB23D1A8867DA25F04B690663C36C1CD1B7D0A8C19CD9F6399E089FE713F5D43C6DD28C179D469897CD29E29A747BCB842F9AFA32D8A82E3F54B7CF0071F3192E047BDF8FF04B6BB1028069CA184AF06D0810DA2C23D8B74C617D6209F89B1737F3FBE565E9D49509C71E0B8FF48FBCB6C1C79B882A0D29E9E0C863865533CF0E105E5AD501B235A499043A4DC29714C503B73CC8A928964ED1E6171E782E0E026BCD270954C06EFE8F45B0C05BFBD0F7E7DCB463353BDB3868AF9670B0C4EA49C59649928FFCA1B81B72048560FEFD6757C7E36278D498B55FB705F679897093CB10BF596227BECA3F2D37CEF13BEF6DA50FFA2058B55A85EFABB94DC7E0E55240F5C14F6CA27751E83C18D35988611905CCD65FDCB1898D602BFBDA78A607580091565255F43A7B6ED6D2E143BBB0EB8632F4CE38E6E497471643A71EE628BA1E5C8E0973E74CFA9B0F46C049D0A3A4D219C0A16125B48F9BCA39A1EED68AB4971BB2E75F820446D456F3EC767F6280B8327DA89BC0D6D043EE8C782D20508EFBBC3FAB515BD64FC25B6137F5F77E274367C13E648671D7C7034336D2C7A2358EE8E3F5A6A5E77971E12F0C989DD386255F40D055DE77DFB2E65139D54731F268F9D5C97DA4868337171DDC6524BE183C187E03B90A2F63B261992D281F908EBD953156B5109EA362F9DA854229404C14795866D6EF8799508BDA1C48E97D129D5F06A670D392957E55F240A480EE8C7DE217A5312DEEC33BA22A48A61DF8553A7E0630B6BD2E2B1F8994C4B3C23B7AD38039413FB790A390BC649FFEB11F1319A503DFFBC10DB723565DC2D17E809F4128F9C53012FB3E5E01F2C37551817C4C654333627CA3CD456A533AF6EEA48280D9F0802E6B785CD9665C9E8E5222779053B17600017932A92830A96FD5A4BAA0811697C812D0FDDB4335DBAF4CF57614C30F9BA945039770B992FF6854A00E410BEB84C9363AA0EE5ABB0398EAEB3C2899FD10E4E6C68C05DFCE03B2BF589647CDC59B891D1012D4F3816FD109763FBC45BFC1EBE7DC07A675A2D9490E9370CA8C0D0F29A881E75AE8F8C0EE6C01A8B917124630222354DCEF430B056BFBCCB36FDCD3B13056CF8BEFE30E3CB8F6EA80A74444DA47E0A760BE3F7F770DD63EF73479E457814FFE5BED8D10CA83121C6EBB18DBA9F2002D543454002FB1BC19FFAE924FD565A69883EE37DB7435DCB4BF6F313427D6ED89834E4AFE1AD2ED92C80245A638D28B9FF03FB2977C847C9E326FD31D44851C4554CA21610496D83585B35FF1D30E24938C75B9431C4254A5B04E94F308734628F419B55D651814A983CED9D1292CEDC762DC908AAD105E0A28867919405B045F85881DC1D6876F1DFF67537B4C7D2B2A67D54E0DD2CBB111DA8BE4D5351310D749254E5556559DB1E963565F2239960C5CAF2D51324E84D4DE74167338598055C676B4E28A88D99426815B57A08F85F1FF1D2EB669D64DFE08D9DD30EAC33245BAF6EEA72A952A8A6596277F4D8CADBBA400376B9E3B4BB41DDF78B4123F2B4E00A8E44D4A2AF13688CCF1B48B6ADD808DEF70151233ED9F4339D21CCCB257574BB3EA2A0D3AAB1516499E8BDA8FEEF0FB44676A977602EBD3F188F54008802658CC447A5BD9C5F45A078C141EC091CC2F12244CD9B0248F2D4604D22F051DA35EBC4C6B5B1D032091411ABB062F31D8C4B8FB5DABDEE3A5389F975EFA563674C39344509955842A70CF2BBD555C2FC5A5FE29667AE036A30DE5C1DF4873F0BDFE701735F5D6D6EE1E753EE181F08BF97FE0D2EA1434E5DBC83A266F44A3A0AEB1ADAEE155AEA677E83E9B5FBBFFDD33550682E821A16BAD516DE49B4EBF2DB9D4F9E05F24E1FF02C9F48B7FE23648ADD5742F715C74A7910CD3C255B06F6B74BE7D9604ACB2A88577DF5DC933788014C3950BB933EB366AFE8D11CD6677E126BDBEF8624B0C42E12E'
				context:   '6E62562D93E29B0DEB2AC27E3FD529ADB52AF8F5A6DA1824CA9790C8121CDEF63FB82CBF730361CF4792D1EC24B1B6B500BEE1571749549A21CA30F5B1E3A0BD16E62FF58A'
				hashalg:   'SHA2-512/224'
				signature: '14C021F9F272E52E01235B92278AB63B1F6E5FBCEE42D6960EDEC79F4899B3246E79167B4AD0458A05890BE0F41E96D71C623417BD9B2079709DADA67582EF44EECC976F3739E44BBAB78297E28A645F356E06095E5305A2905FE04840D6DD3E773B7BE0FB8AE34DFACCF4F2B0C2018A6606B442AE12BC36A432E8E24B50F3DA30874C48DDCF73C41AE9DCE0C1A4D36CA215754665FCB049D2230C2B7B9B643D75113364F3C3CB89AFFC6DA545FB228971FD06D2CF69A06010BC0E6887A643FDD68BB6F5558F5FE4485A8F4F475CF25B38D828E3BDC8855696F5717476AA9AF3011A4043B25AFF1B5B4660533A98A445C98D164F987EB4E2621515AE04291857BC029113EA0CF0D7C0CF07C58440E676CD7963EBB0C69A720861C7568885E6EFF70AA89FCF8190E0FD8EB0765D11A1391182CE96A42D65CA772F6E639FC7D317B1B8998F3F9F93E51B45E6AAD70542DA3E5F6668D97CC377EF49B79A525A3C06260A8AD93E5E2E35E90B664B3A7F6518BAA44613AC1F760AF83494DCA838ADF1AAB1308B884556749749930B4B23B11DFAE60CAA09A4FBDBEEE735B1A56FC0DCAF41840AF804EFC12F58B2853731CE62066F2877D454595AC18E267EA722D09B3302BD1045237B8EF3697E969D77F8695516E1B186EEB2FF4EDE19CE95887F5F9F2F0A4AFDBADAA76F6257040C421CD8CB3984CDD7F067589013556161DF0322A75D08E15D9FF271F9FDEA45526F55E14F3298843EACED3691412B63FC8A7C131BF40CBBB7ACB384B187309262783B46E614329F2E877A9C090D0B415B9E221A64871646D41B4F9BA86AE9D71F48C57286E26057FC7FB717ABBE882A4424B2BCE4280E2B60E0067D5B5DA945EB102242E697536AAEAC53DB667D878B02E29A19D31A3B46287DE4A755FAE6B87E49B29600C285F55F3D402093F95D0D20B7F832DE90AD4DB14BFFE0A42ACA391567C02A679358387926F7BF1D54FA7BC05AE2B99F409ECE732562FE794CF5F5C65C2C97B13B565A6E95763534B34D9F2A8ABBE2CC463777A80890E94DC0AF9DCB9349D98183D2648D8F4694E61ADD944F12919EF6E6B0D0A9D431FAFA216AEC8FA31EB8EC9FCBCD1C1B5BB6225EDE094AC81FA6CCA0C534365C268D69BB01A9BFE186D2DB6BA7F40C182F8BC2698FD81E05C315C743C1EC2E3606E2D750430BEF526153D38EFCCA40FC095281B8A08A8A509D433909FF2E8505DD95387DE275B412E4B00C3773D7BC98714394C2FD3939575AB55D463844EB4E133C4CEE387A142D10AA97A6967304E5B34B6FF64EF0DE9DBA6D860F22EDC9A35DDF56359C4578DBFF2EAE42B46EC228D6703992E5CA9C07A3BAD255F0A05FADF719A9B6CCA6F32338E19D4D55B410AC2194D347E1A6987072053209DC9513CAB714A7DF672378997AE2A09AAE31AABE2044CCD978433E2D1B16EB34B0780BAF976564C8DD4C1C2A74C56CB498EB35C9906F3F9F183AE4D974FDC55F810E280111B1FE3573247B4DA677A06F9D9134FA69619DEBAA0D8481D40EE18E2D215E80A88966E2E0C9B535293A5DEFB3016ED181B4C1C7E32160B428FE065E735E430FDE9D6B2CAED9A42FDB289452ABE029122F0E97B3F2636873B734A18EDC590F27FFA0882B1B4611804569BB93C63A985520B111EB17C73635424AF7DAC99153E75BC57F1AF72527D0860BBAE9F678CD6BE999D671AAEECF13A5E4727997B6191451AF25118E4E6C8D362DF98060487E07302608694309F7CD530DDB32D47BF7191CADE99427902940EEBBC4E6CE361E8BFDEBEDA492B03AA84C72676F0B85B30B13EC9711DDF6687AD75C4B40E683D61713E6B266BCA9E8A9CD45AE90D9C177D89883CE0E17D034D95FF3E711C1A7F5CE8CA7DFEF97D6833047F5C64272476CBDB40922590170456CA16DB04447CB82959527D884575E49DB0607C1FD1E29A5DBBEDA241139FF4CEAB60B1F9BC5E613CB5BB0A837E3034500F3D6226F3AAC348C0B275C5B72F7ED0F2C61B3D45C6DC9135706B516BE7018D8C412FB5E5EBA059FD308436300838420821478E22634ADAA0F8F1A7A29C9C85741C13CD2C8D9F4EEC9BD7BA1A6B1CF25C38ADD692B42095C350B2114DDEDF246139EAAF29ABCAC721DD286B78D56D44C4A9A5CB2EA2166BD7F6D12AD94DFE94A409754BE0E22B59FBE7076BCFCBA8A94AAE0364A72DF86DECD7C42FDCF7DE23C0286631EC6E27AD07E8AB1A8B79DBEADA32386600E1A29D9F27E4F679AF59C6758C36599AFDD09B8D2288D7BAD082781B6A534DFA93206F38E536D30C147F0937E0518D66383A4B4BAEE2CE3680CB3C87AE7ED576E7A7F4E3EEE51A3A482931A7C5EC48A452881046EC24E5E33F56C36B3795C359158824BB13EF59763F21D008FE8698D7EB84BBD354103A8A618349FAA1CCA5CB72B02B93E72369052BC0879F44A725FB30D7D4C99BAF445A9FB10BDCE10DAE653E08F25E527EE849D7CC64822421DF7B5917566C0EEBF1FA45088833BD5622178EB341C7DBEB0A7205BBC9B7E6D4A9D56F445183DBF9A3AFF1D998D1E34DE1892DD7FD1AE548939C31108361912B1600C4DBB545D9CD45BD83B662DA0A16FAB3C0C3FAF138CBE6010F24ACFB1DBB8FD840A840581DBAEBCE0BF3F3F99B88DAB5E84ECFE933E5E21FD79CCC15965F57BDC2280678DC6CC10A615B1B301E8AF25DADB5FFFC80DBCCE13EAA1FC6363CCD6FDB5579F7BDC65D0FB706B384E4E5C815C6D7DD64D15EB95894668DF05DBA68EA0610A1F5ADD4387DFEFAC057787CE01953B15E22FF98B4526382E3B4603BB65B005705ED557F48F77C9545A604BBDCE463582DDB2C1D5806F0A5B89609B530E030E4FA0F7D5E2C1D7BBF8E375F1FAE20E6FC271EC93B6D466FFEAF81435CCFE0EE3751A16A70429939F973E0661F6D66CCA173121058893A92320CA50E07B995FE88127B3DA2EB780DFB2B5498491B89A22B61717449700A098C52169CF176A0E40567E25B3C5C64E95D6AD0C4EC07C861D4E4EC7255741EBAB470D78E73D66FC94CE04497F3B00BF3D8EF4991A9DFD2023DE449C90E6BC3E07892241CA80EFFD16977FBD8B9C1C0BBF2A1170F5E881267DC560A9C995C71DDB4FD3E27BD741594A25F80C705BFCE5143F6A9AE5EF2422AE34AA82D590F7F55631ADEB5B4CAC5228964E797F9400C8454853E55E2ABA9D29430647CA3AB62E27330DD73FC36EF75FA74FCF1FFB40B1C75D0754940CF2E8FD2076242D6F567AD3C80B585C674E375B678414CF19A79BAC4E214B51C6D96DA86B3A5C3B085EE31D1ACD6E64854E79D2459871C4CAFE3054CF390A4BC9CBE5ECC4A1AE8CBA1C58B59A72AF38EF20522BEA92C002EE0B3C07B4FDD9EC48B6CC1897ABE46EA7BBD2202E6FF7C94B432E40230C3CFF2982D684004D027255037EE778B09038A745B390331AAC570666EDFAD8616B9920D8FF13563FCC2C0D1C2A1A274330A6E81086606CDFD291EB03ADFF17F6427C2E24D38158E10185B96ABCB327033FFCCC2F2F1E79BBD6B741F4C4EFF9ABD2F220D5BDD20FFCA070B6981AA408964954F11B69122C9E3DA2A364BBDF079E9A9597BA90C49D31C91BA4EFBEF0366719883508890E9575489ACF508207513FCCA70DEA7BA3AD5BBF390A79ECA87D10A8E425C5E9629A79EDBF4471FAF78295594FF570BC668A98B2CC6395C121B5E45B940AAD28D7244EB4F4F8FCE59E0EFE72A71B04CD11E990C641E7C44340DFA770ED30264A435F2C17326777753A9FABBF32CF592BBB69C2A24ED5CB056E9A93CC5EFCF37CEA3D407E4531C0CEAB810ED06BF244AC19B9CE3DD9264A013E12A52BE4DDCE33F1879EB5DE81E7E95ADE4C795DBF051FF0120802D3B5401F9B20B062E9A01FBFD387F8265F0852BFB703929B7926873D3EEFAFD24104E59F83E630F6882A9DB798440F99DD134524B4A5F04ED1A78CEF15BF3C5E65ADBC1221C33FA33E2851FE8671B6DA3C909CA66B8204AD5165CA2EB1C92386D6ED63E6722FA8D7BAEE3411C206B9391FFB31F4C079B2D243396347A185B208D933E9E3E509206E9460808ECF4F0D35C6C08110FF872577DD8082B031D62C2F98501482360A30E0C3A761BFF99D4BA131365DAC9C67F8D72F6B6562F3EAE00016E044344A6C4236B194DAB5FF87E8E2E76918795823016962368594A20D116399FCD1AE8B4774BA55503C1D0EE8FCDA3EA1596FFC58F1E15B998BD619610CE9224EB8005BF28375EC0B6F18759D272400876AD3983D29DC00A9DBE455942D40A7B3F87BDD16A0D889A84B49265331F667AEA5109BCDE60AFDE19E8BEFBD789DFFB941FF078B482B49C6A42822B0703DFC7B7C910D203B4314B361123457D454571C01B582A26989C5D9186A68ABAE6E24C4C4D902767BCC0BD124657F58B26F12A3E5FAFF3035C8AA6E511573337E8608EE100A1676D098EBC5E39ACD701626B04D317C53C53321F1BFA000D20F75824A2E9789D9F1B81D64E1D27088E00E09EEB4EE128AEA01ADAE8AFA045E02F24466E7115E6C9760CAC177640824E35F69254DCA2B2BA9AA90C580FB87F1382100732D7EAB0B5D70260AC30A4984401FEB47C30CE57A49B6828AE0D04B57CCDEE221B5E3D433C1A6C92516FE92E2234D12749FB6B939364EE1533745E5C32CC88FCC6B322E0CDFA280E689391E0F81A3D5BA56BFF8F724D147676E5B08124D24639814DF103454E8B07A49D4C97258B8E078F677D2CE2C1312EABED6DED2DE3CECF1D12A12EF8A4C27FBDD7DE0F0E345AD4F5E7A2C82E605DA53E90BC045AB5EE6C749031732B644A6E4EEAB5AD1145C111EF7BE3370FDE0EF5EF29FC5226BF5C18318167E092847583CFED623BC90016B4F7ED64474A517E2545A24924B42922FF042C37112DDB6371A319394C628F354C12DEAE0527BAD6D6D6B9130D80CF8EC485654B3665CB5717FA4D4BBC55CFE6B570CF1406D926C3541641A0FE6527624013EDC7149D4C4FF8CFD15D180D15AFFA9522355086F0252B6466012C1251738AE239EE17DC8B1893DB3EB698376CB1B1B1EE00FC42A7DAA4011D2A272C966F154BB9CC910227A9422FB53BFB310CD652F1E65C1DA2BE2C9142FF68A4968E65D430C62B85F2A5932EF61B768CF15F334F7B0046E47F03A6920709EF7271C6D146CA25E5465EBD3AEA77FFB090D69642D251337B91906E2009A8542686B047DE8BA9B156FC51CF3C5108F8FC6AFB94D6D9F8C42CA7F7962D8D16F16548FF68BAC23038CAD3737FE37E0F08BBAB38465FBAEDE4161C21DCF359EBEBBD73D5B26317F5753657FB9C615B16B9F86CDCF9BB1FFBC5775DB2B19B053EEA4D9F83EFAA1A6FB6A86042AD393832FDCA4736B678CF34D7110174670C68E6EA71B4CFFEAE38F0C967F6181C34B2CFA6BA7FC11ED3D312BB0B8B9E6BCE0DB81589314B48B5145C3EBE9A2F2E02808EF7BD0084DA7995429B9782F6020D07D7F40F262B7FC38EA5D222D548566451EC2BD721130590EFB24947F3E8678AFEB2F574D7036F3CE4A64A44256BF0276AA00BD859B56FE7B494D04FAB0E1EDFE9BCAC06B77E31D0A28CB3447B94B25196D71B045DE1F5A91071585211164993737087531CB864B216C6466C6C51C1D87C25E14F247C5FC413F323E6326A6371D3D9FBD5DEAF09F4690D77755A5CC432BF30B556E084095F2038E00C634F27A906C4C78BDD6A44E566B6BD00978BA34322386051204E4BFC78C29DCF2197650CCB54DE33A66B658F8467488C7B65AB1DD23441ECAA3A578F8299DE0F1CC1DB44B101819CAA29B7A475BDA72D3F3544FA39D12DCC73D936BBBED8350D9A915F454E850416984A06EF3A02AFA322D4E1BECACE789CC9DC04B62B183CFEC2D202A436CF14E76E41A19762755C5A5092E63D7E42F0754A5D5C6F5EDC4987A4E4DBBBBF2196D84EED6E7D06F24C4642171EC7E9BB87AD27C971C48C9017D89E18D4160D46589E381C61231D4B460160D2D70557281A04A9B9DAEFEC0E89E792D58C298DECB78F1AF270AEE9F17F26C9AC30B722D1C5FA866BEB9B8ABEF234A5D27A44B141E6C82AE47F0088080174C00687B9074E4AECD99EA0374DAE543068FB68271307565EF108B08F9B66286C08E6DEA4681E59DD6C993E8B08E4B97818AAFC6207AEDDB037A045F96E8348DBA2E2E075FB0CEE536E32647782FC3E17897F105E6682A600124453BB58EF061FC7704476057B7B3E7D27F54093EC4AA5120166ABD61DCAF61859988AA24F69E8FFEEB591CF07ABB223F2702F6534B74B9FCF51D5055DE317DE3D82BDAEAFC2E5D4D851A25F20C39293F69EC0B344E7CBF56A44C7980C2966B065B267E20AA27B4AD0C2BB9369AAB192F30B0B3CBF9354BE4D9134E95C3A15754036D420E0AC466E9A470152574B03C4C60AA94D47D9D22934C9D136E4DAC9CCF6D1219691B219A34779C0C2E4BDDF4273C135B82A96BF942D53DAC61C28D4FCFFE2D7961B3959A045673E65D08982A0161CEFDEF1F9F182CF7E3B4B477A3DA9C426A0276601F68A1265A24F575BF982BAE922773DBA1CEEA4444563C09E1CF959B97755D17BDA4FE95E063DBA1AC8C9E5F7DD6AF3B84E0F6211788D1185D7DE72B899FAAED72871BE7719FC1A17299EA38829547F7882E448F43E3AC7DB22D9BA182FEC5CF9C2231506C06DAEAFBD5E8E35F695B024AD6EC52FDF429E21A2D0CC8A1BC6B8C9180F9D81B95109FEFB0631916CEA0B6BAD2B9C6630F55C85A88F8F6DCBF57B997D56CF490031ECE4CFB8E7B95E16814414AE15B3FA74C0AAC117766CA6263C43E62C5BAB08A4E96E901597406509B899DBF065FD076FC0290F909BE89B8CD0B95B795600E9B796985A254BA6454552B0564348264F9E3A64806E33D9B1036D4404CBB2D4FB1FFA8DBF7F687B402880548BECD22A2DAC17AE6E8D121BD4B387FB763607E2D419FC3D88A1CAA3E194C43F0E54EF9ED038A572D0A414A556E84114BFB5A2FA5DE02852A0253ED8DB190FF4445B845BDCCA9E4197A4DE32743FCEC16516194F7CAE99800E17AEAD3D6ADB00B8480A9622C1ADC1A47DCDB7689B9100CB2E9695FF4E7B1690C30746C53444997603D9BF10AFCC5E4063F4722CED53822C827A9AB45F4980D2CF14DD32C70E2311F58FDB4FD20437F9C4A090C0EFFED00F881A39C2C435EE583B31AFB975A27C2F30135314FAAE1AA2F3A20BEE13EE8572DDC52AF7005B1CD8C1571B7857ACD6246EB7D4E1DB6C001F69DEDACFC34E0B9F6D4A765992EF1C9518A2AA6BEA0CC06B533CD4D9D6D59FEFE8961B8D3C86B5CA2F23AB7D42EAAF9E3F0823274127D93FC7541970EB3F1D871F6C88D4A2DAD5CCCE0B008B6B3BCDEE18ADE6E1B7A237BA7FBCE867C680EE45593A337C258F937DCF5CF4BE0BEE09BF5F641BADA5351FE76439E9971F708FAEC7F6332F20815563B0F29E4F0B7684DBFC417AC53B7EE98A88BE5AD335F8D1D737FBA3EE6CD4D8C615F5C0A294EE6CC82D7EBDC1264E714F612614AD6EAA3237170363CC15B6D614A42346E91C71EFE436CD51818743CCD3B719BCBC0B2CB8E51AB60FE9ABCCE422D43EE0AC496F3DD86427CDA5B7383CECCBF663F4736A12863CFE2B5C262632C583A453B9219EFCB12051AEE36B279F9353B099EBEC568D40E65713465587914D62AE8B350C244B19E94610F88211AE11C77A164DAD2B0D2EC3516F8E93C22D77E1507D24D2B6005B58D0A71A4FAA7A2853B2FDA250F3BC8B8CEE4966416C1D5E0A99926A9293CBDA078A0B3D361386DFA7694115069CB482C49154DCBAC42EBCC46958A08778FEDC934724BAB010E6FE1FD9E16F95933936017A7303F32461D1AC5DC09082863CF0D91E249E0128B6194805E8F6BBF874F3FD07B424B4D5EB5340128E39D15C0378914E435AB31BA90E2ED7E15F510892CF6EFDA308126FBF716AC38001D41C74EB4F25A42A0A0155E2B713AEC108AB773809C11D88C957B71BC1A2E6E77296C91FAD9EA003ABFC96E00C87BFC16E6E6D1A3B5758A754B2206F782C1F5BA3C2952BC1E131DF069A8ACACD552A563BA78FAC0F71D9FC22CE8AC3D44ADC2ABF60F985BDCAA21D815049B053B625BE1CB06D8952182BDE9960CB225DAB4B6C8A772D4239AB89359E2170AB459D014454B0E204CFD14EF5E242F20CC397C495B2A54DF7B4969148446B971CF22A5D67C9B0F3D6862A1D3853040AB141875F6D63186641CE279D1837D7815E4FF565FA96EEC3BF5833A2C7C8B3BA023991396672949984AD89548ED580C5274B7BEEAFD2296E4A5C13A757C5AA937C8A915C49496731E6299CEE764862B60B5C18D37FBD3E3680735F1E947D8CB5C9AC3C97850DD77C7F33943DB844A5AC50CF0941FF0B78DC464E8D3A0A702660B9F13B22E7A219DF53893392176F1A857900BEB0C748D02F546DBAE6B6E870E7845F4BE3303F382E14C6A6CC06B15CF1FA3F69DAA2CDE0BA282CFF1D90B5DDC0F179C8530945DE4C34039C1EAFDF8C4832D85DAFDE85095CBD2082EF2B72685051C323BDBC3E7A821183C85AD349196EEC727C057FFF991A8A1931520486D8DD8052E6E8E30CC1A7F04FE31CB39BA909976D9ED91CD7281BABBEA006D28DCFDD29C9A119E8E0BEF24B7A72C60724F61B4EEDAFA70B3CF34371E01FC18FA7EDE8F5E48A4F065A542228646466E7DAF5560BE06131D2DB78AA3A7042166F3596745C2B0706646E138BC5D5D61FDB388E06DB06E05CAB7900283B2B9B3BC69FBAADEAAC6B91381734F62F4952F62F06BD21C15C2C0743AA85634C0369BDF75F6FA6B57607A34D25D4F58F425F974E85E81776247256487A36A21A817F84A82DD4DD1C323137A374C871F3BE82E6B699DD9BFBB4BE2472F5A9DD013D02EAB06FEDC655A339A88CA5F2568074E5E874B5CE3E5BD3EEFC4273878D5C21E0D44AB8D6684B74FFF7BAD71BBC7FA78118780ADC184D3EBC51D0BDB26065DB9CE81E7EC369462A6806272D773E654A46C2ABEDD470A3B52D2DC591BCEA42A32E2B9948C53B182CD235DA339634FB95DD73F097E1744CEE2D1476DFAAF5B2F82CC438F927DB8D27DA4B02A98BB7FAB8C867B5A1008BA8CAC18B3847D6335A7ACAF4A0B8322D33117B66ADAA2127ACE4E98C21C13EC75FFF807241AD84C6CFE2492223ADEDB9C804C22E7532CAA4D63DB7A4CBD4E5F6C45B7B8CAF4C1322FDB32FD08F8D055F4A2055FA203C9C4D95457CA7855ED7F282E6E207E7AD36BCB86F4484FD700742E641CBA9DC03A2E6A4402B05B498175F4BD6F2D5D9A25D0D88DC1416DB0C927E266747273822CDD1CF50B62E9613E458F927838091AC75A2A0BC01A8676C9601F8B476B8C46F6865F0B4D5B81694EA3602A23F1167278EC56B551A3784909C9E5AA5A82196C3A9C91398865DAFCBB2DC0F58DD2A093CD4F8F3EED13176336CD854B4D766B505FAD90BCCD5FA3BE8A87617FC49191F3D7656CF4FC431EDEFE241A43990ADB37A78D55498EAADF705A1F0D8AEF204162B4E8E979D82459A1FAE9EC091CCECCD98D14D1A32D3C1D45B24A13D56D4D35230D3F94F78D8149243856D3AA733879D11E7AF840D946E1117C840F97DDD2564C63B4EBBFAB4C55C4D6AE6608203310F88AF7A9A28999C923FB1291A54C374486AC97C6727A5875AEDDD867080EC417930D061C5A4208B52DB2ED22E05429EE86862F98D0F710803F043E98FA31370795B13893BF342C92CF5915EFFD5245DCBC7DBB8A1C57607220A4EE993E67CDC88418A76D127B6399FE6D457DCBA140DB4F117CC49444512F3D5ADE21EF1D026DFB021A7D8592E073D8DB43538294D2E293CEB61583E1ABA0B863C358E707E5A9B689FC19C741E454B0741B86F07F64D6659D11ECEF5B451BC80C5156236980AE0BD7027F657537B9AE051A623DCA7A26753B8B8C7789C0FEAC3BA2830D2803DB8357A643E1F833DD4FC105C72CC19AEB3DB422268C792205386D34A777C3485CECD4F08494B846BE597BA3DB8F1D64E4D8D14A58A2BAEA481A82D6F3BD193F2283DA970BC81A37757E77912C676BB241EBD769080123EB69840A980EB80D4BA35FEE05C41EA04AAF3969266583173A496D6198DE389EF6E149DF13AE6E20CA9EC6C42355E75A6F88459CA3F63835F073B3FCA57E67CAC41BBAA12CD97218D35251A2CCB5AA4F7826EB57063502F9B61297A65AD6BDE642054C3C4B429DF1CD6060A2B6E1338EC6F30BC52855168AE7AA8879AE71B1BB9A56D3E7615FC53CB3112F92643AAFFE59873532A41C93A7C8008AFF21DF69B5314B97917CBFE1BBCC02D9994B8EB85CCD28ADB17231874576CAD4A6F3B95B15D80AADE8CA63C6136824CB9E289B62833AA5BAE7C74BF79FAD2C37998499A16DE4B7F7C66A7800B66F3536DD7F4EE28D22700BD260720F509A09753B0DAC8FD89D652717B71147B14D7EF3B3E5BD4E15008AC949EE3A75ECA555441E66B5BE149A65F3BEFA795A5824AB9975D671E078D355EDF77726D824F1A08AD39E1FC8F22AB2B595661962238B73E386878DE10FA8EEAEE9813078272EBBD117264759E7734017DA7118E3B99ADE984C3BD540467A94E2138F2593E10C724F8FCEC6183F73F491FC3775B96CBBB7A3AFB08AD328F4E0809B12717FFD1228658ED013E86C90BE320F2A044C83F09D13683D47B4F0E6A90A5372714A103A3B4846C444B5CC4C933DA2885C7BC505E35F72559CE68439AFD2993D67C6C7BD7C2151964628EE4C6D471D91047B3BE2AFCBD841D939BC9EAEAF2E163309A2D79E1AE9B22F3C4B2556270A73FC9A6E14991C66024B744660AB92D55F8EDF282CAE85054AC180E455E2CDE77C9E70984242F3639B3C404824BD3CFA88F3CB62AE1EF3BF3A76267AF409B0D870EB022AE7EFD2DB3030368956C2E716AB24D1EC2B94F8A6F71ACA82638F98DEA3D8587FCB1646294A2594C7EB3BAA3695B2B91C48472735010DE769B6D363FE816B5D9624468F3343D4804E5F3C53405091845F53470DC1EFE91BAC62DECBB92C8CDA81A3A4D295743AADCE8546B1EB5222B23E4F8D6E67BDE334A0E934937AF5ABF6E587F7C852FA8A904DA46E55F67E1ACBE900B2DB67E3D8D3E279D57F6CF0105FE2CA0F9B5FA345366E954E172916E2AFF7B75CBC57EAB537657F089A717C02B5D25B65A96DA70AA0587A08F7B7DE279B5D4CE81E54ED9F9DA502238EB874159E85C5331F6609A43F79D8D5918425FD7A19F2417BF98B344837B918F130E052EA537BEAA95D61A414F628113C80DC66C84BB96306BD1E8D0ED46FCA51F02DD2F1464573D134BA93B6ADD8F54274E3A6A0319C29924FAF23F1F2FD25BECFCFFB9BB78D47BE200183F5D31D8224CA88C1C4592C03A0817113C412E6D5C0F7A3B42689886C56C5F0D594C30DD498839C462C04D199A4503C5BCD70067FE7A900A24BE0569CBA9848AFE4D1DFB91FB0E004A5FF74D1E43D291DDC0E631BC1E093FF16D44A60468D7D174BD0ACFE34CC868AB1C5932DCE40251BFD4096BEF35A7F65A35A686F699104F1C57EC2790DA0B8835A60C398A1BE37E6661592D11C347BE83F39D77295B2288388F089C13E5094D1EA70A77161D52AD190E0DBBBFD8A2E6D250EB03654A50F240AACEC785EB91E92557EA0B5439B9AA1401DE498C385CF2A1CBC5E8493A24DA552B5C36DF9F9A13E0A659EE73159AC68BC18376B56EDBB7BB732976342AC4D30FE5A94F7739272F35166E1AD70A83BCF30AC4047679036F631D2A75E60F7B0453620C6E121E04E31C859246AAC3C990E0D7BF9DE7F758BEFF80F57174B306FF7DEE47412A22B3D1BB131EFC3B336CF984401691E41045D2560AF1887E790A4631AD8CA8C51879BB1C67D34FD6C1855880571FC5BEE634E8AEA0E0A284BC16C20F7444466E374A6729C3B4AE0AC4E645603EB54DB5A7AF6A9D6F5B19D61AA2E871EF029E0825C7B9171F1EFCD4374C768853053E0914F8649485D205C70E39DDBB6BB88C153A8CBD480B1A0207D29DD63265EC17D2C709040B158E0B97796BDB995D1A7BDF91E7E14BA89B88FF72D4C90A18CB802ED9A73234148C74C89E9DC3E4A42102ED9411B9F7578D3EE20F13385A4D3C1C75BECE42A558668D5E73F94DB51A9560545159BF35D9DCB1C23BE4D78E5E97A48D5AB8335C35F33E00FA3E2750D3D862FD09A5F6776B84666394B63FCF3C28DDE27046E1E66DAF38A6D88B59B7446530ED46A8DFCAAEFB0128262F0CC030CA55167CA35B535F14A4BC097CD91CBC65371F8A6D6ED2297EFDEE6774782441DA726CC80AA79045F6E268361019A0B76627B61C7773D6A53208EFB4A64986AB46F5A93A25B780A3926F23AB961983B4D79AC1C928C11C33EFE7F4B0E79286D5BAF5E37C9A1C64717C43736779AFB77FF9830ADE8D2480A158D39587795287C440943707F95B9ED4038168D22C32F7096870BDB61ADDE6D83449DFDDFA382005B1F503D1DD23290771371B67F1BCBDF0AD5B75B1FD899F71932B2D8C84603F9D3AAC4CDA74ACE0F91208FF25891EA151EB1121C14688390352305A283466F6BCE7EF741E6719456C911C86DCBD9523D1AED3228583A80FF1C8BB619AB6DFDF49B47F1B3EDBB16B7A8DAE3E2A5B63D7B4B0BFAC069653ED30855184B5F1E86CC0813C4E75B4FD5402E6AA470E989B3937E5F26E23F5F025EBAABC9AA3504E6F566A02F05249F2C4981B780386A2C5F92C61A4077F99E95E2A794AC88C30B06D27D30A2D9E62359D6791C821D82D3B9E8ECE6BAEC4F6EB07CD0FD4F913EA48923ACCB4219DAF972172A8EA9FD91C3EB440CD42B228B0ACC78D0D889707568F32D33604EE3F49DFD1EEE68D76119A0B79317803F01309A6D8DB7E7FDA8735AB8F640B0E4B37E4A2D29B800E24CE31183F87C5458E9F69EDD24D66CE12578641073DCA0D3F2333EC42FFB4684735A6FA8DC0E7F9C1EC06E35C69C4BE4C6112305FD0C0596258E416E55B76E95C3E92BF7171A42AF1DED0823E905A244FF0F8CF6357D2A3591EDAA197BAA16516A63154FB27DF01DE255A156ED8F2A00ABED9B0B42318BC1C2BB27A1D9BAB2CC185BDA3679548D43F7B6EDE90E4F5CC1433F785E64814AAE7439613B504DDE4B643C1BF91E8439C3DF0A7F971B9D534EEE36A7D0D6AB65A9EEA8A668AFDA15D0DC18F029B8EB5F935E31D10B4C8AD7F14C2FCC8E1E6BCE3B927F04EE3F8C16C36F945F9DC110A881FEBEB3BE7FE53648A52CB36BF88ABAD7855186D5A0C37B12FECDB38A4682ABF1B2AD753DADE7AE51EFA98D5D2CC890E9CA901D8D0DDA1ECFD0165A9B946ECA5DA79ACB96E565EEF8C92ECC56B0296AAFFCAA79311525817654085E609D5AB7E895148635BBBC18B90E5DE5FB7C85505D124089E0DC644F7849D7DB5CF46FDC87FD7D77676A38343E5A2EBB2BF5BE481095065E38A18D8E949A1CAB5B25FE9725BA26EC09E5809858CA3A1CA7A842DC63784AFC6CDEBEB94F76CA9DB31C87229531D8B4B148E7114229073D014BB98F16ED473637BDB23EA0AB8009DEBEAE8F189F2F933C321B86EADA968C4217C22B7B4A71964477E20E878E71DEC1C8A1F9217B067CF16A59CBA6BCF014F04A9BB3151AB9E3436194763C24A44E36D47FE78921FD16F7D703C39BE1F2E4BC962B57AD7C9ADD81DC5FF64B014337F71BEEED68A03B997B6449DE22BB6FC2956F38F1A72865655EABD402E52E706867FD147106A90CF84005DC0F430D976E1253823C9489B54E4FB876A831B58D34921DFB21CE643278CA7FF43FD2B4711E19E27B1D6FFF91D3012D604F6828B7C5066FA93F933447C9904037C1F45C774275341DB4199498AB145862CBB4C7D8B1DBB05448DFEE2F5B261F54CFAB52AF1A4A926111BCB8A2CFD6B9731EBC8C9E408128D045881F212A68E06D39279717DDDFD8D5D2317B4348C8741734EC8C6DE929D4751F13EC9A3F58E210F51F69CEC6C13F6ABDFB6BA09DB9DA11FE7B9E6456EA2A41CA10FAB46C90E3A77928475DD922237E32A5163876BFB539F09B6AF6CD6D8D183CA24FAD700EE8D6741B3DE93D4919035151B3493C64BD23F920BB195D2C4F5220B3F5781A1293117199280B5EC08F96969045F1A609E5D25BDEE21918A62318895F1F49F6B58AD9030B6456C9802DDCADFDA1978020D0D8AF3E5376DC4ECF0F6C6AD155D8BE0B0B05616101B94C38EB644D32858855DB9DCB9F6B5A9048267585978EEFFE93702D82C54259BE3BBEDCED25EE25CB6C94CE5800D3BA4708E104F666455C984B3AF94E9AF0DEFBED1409B23679E7C78A82D69847B2231D0FA53DF78036176976F5953140239F7C97684B893E684C5F7402FCFF6DAE3189EAAC34F7D3BB437577F76DD2824099E8509A12B04F48B209BA1DA1ADE6DDF2AD3B3DAF0C17A9245FE6A2E5D900245A29485122F114810CCD15AA7A7D029691A6A3AF7CB81B93DC21853B5C4F2711D0BFA187E5C1044745299827F6C9D8F31AA9BDF414B93EDECB9D87D161F994ED176945C3F67B1F7D5DBC03C778BAF0E56549590F88C05E459B6AD591132B27BE97148ED898EBB280CDD903F727F49CF048A04F1A1AC4E1D9A789A5264DC34304081083534781A7E2209FD12156474E9CBAF8970F7752882D29C16B91888C38E5F5038E522E4C38385F4267AF23CFD3E16343A034460C60DC6A573AAD1DB3A580291CFE202E2DF23E135CDD119475EDFCB22566FBB9317FA1A1D13D6F956EAFFDFE79EDB102502A7474E79053E6A446B59B7400575518861DA3FC7D10DB98778E8EDD11E4F355D6587303656833C60C1E1DEA6A61401BDE8012D285B55455ECD5954EDF0A29F32C5ED2FFEC7C60F57800B4EA7841A9187567AD0CC2A6D2E95E177C26347E8FCECA3D50B7837AFCF0D961EEACEC0B38ECE51B5F77A03F117D7087AFDF12D4E48F57791DDEFC1DC136DB167B20672BDACD61D2284EDF62E7185F806B4652106E272D0C472E7BA053504472E8932C2499AF6DB3955B3480885CD2A3184FA2B2FA817843B956B36AA95AE586D8CB9CAF8B8F98AAD9C01870F7E898808FD1610E1063BB2A9476A13ECE915BB0849819516686AFB7B8FBEB0AF075F5113B671D8BE445F32BB8A36352A38C2734647A2C02F3EA3CA132400412CFAE9A2CF8110EBD442B56BB4BAB6352F0A419CEA3B088232F24513D16725AE5B6A894C9947E6F7987F9B97BBF776DB26141FBE2A4B57DE9F6F85E9A88871020C70B7A509E6D53AC75158500CE5587E58CC48880A47895F4E55934332FDCFB312FC300CEC2CEB3D7E83E34BCC75FBAEB8DB1A014A90DA3EDB450BA37FC29EC248DF0E8509AE2B81C7DA7319187D645E369637959C50A24E2DE230C2F0435F7464C1E1598332542526DB7BEEEA4DF096B9CD4E29F02DB37E3EFDAFF194DBDA62BD19A383A88D234F75BA7CED8D8B5F1230BFD61569FB730396383C70081295A8024F91B388A99DECB5DCA36EE1B413C6F2279EE747758DE555F9448E7C8C879C4AB03107D1AC60E7C11CDE9866F09CB9ABA4441156485FB5AB98B7D8A85CE64E77BDB483E5C2288D1A429AC23D6A93C914416547AD896AC94AEEEA16E2C41D2B6228DDAAD73E6C313FBE8EBF11E9DB5893EA058900BD22A4EA7B3612E2D1091A264C48FB96E96A131EF463EAD235DDF3E06F472B894B0C812B8538C681104CA2C38FE4207B1F96D4262FE836E3FF1AFAF82FC63392A3F313C0619AC56C3A8D28C723534B7C3382BC736583641001E70A0AC2C01409F902ABF53D435BD11E3318832CDE4387A8C89499BA51291CF7B94E00751B9B0F7EE2E7DEB6BADBC7828727829107F56BC2563ACC948BB622426059163C41B17392A00630BA040A495EE8AF7CF39704F99C71985198B5AB269BA026DE744D1AB9AF6D4726283F6E830C52158E8751547C913B3ED33903CA5903A2EDBF81CC2B9C218163DF75B117727C20D8738934650D9B754265D3E3831FA88D6A91DBC42F4B5C0755D03A8A7D654037605D9D12183154A73D3FCE2AC47ABAE488EDE78567CF7633DBE4CFEF352FC62E31FA51F1464551F494A51B0F0B5413863343441C3ECF7FD7D50DA3B3F174B4451783A0C20F1133ABC57A547A79C9630F5EC79EC5C0041EFB6093FC78B9AE2116CDCAF92E0ABF3126439A89154BB459E37A866801F0DC3590BEC7A3D792BED28B59D483F0C0E13B2C098E9133C4AA709C84E59C5B122F52CDBD838056E3F601007FD855B9312C4F7A59E583E35644FAD767FBF7077C4F1285A13EAA2C7217BC1951363934867C3B072518416004D1CC78EACFAFE3689076F95963B12C09842665114F75CB1D05A16C07D984A810AC88931838EA24D26958FB1523AD2927F9EBA57E2DF15943D60EBD00902C2988E09E8ED4EAF5D3125199060899A217DCEBA163717F89C553BD578888DFA0CC7652353DFFB676840565AD18DA5AEEE2301896F3BF5679B17FEC3303423A237AF797784ADD1644EC5636961B20951AFDD439649F8157A10D94CBDC9EEDC0BC8EE4E97D45F9BFE486778E4119111145B3D22EBD0F0326F97658756AFDC7E170B8091995578FCB2110397F04B2758409A9D8280A60375129804CEBB2BA1A467B5E0D4E24E7BF8E0DD4D91CA34A86E4327D11B2B40066B596D3DC9B6322535B4C8BA3B2AD03D29E455828664F3C055D7E957CBB5C47C7B7E475476A01B45BE7DF537AC29767A361821F59DDA64F68F1660A7652C1B860963E6D0C17BD52CEB2B53ADC856FF6AAC97DD16C1376A51A667177156775DDC900610A8F8F59B9EF7705CD486C069F59E29B239B1307E9CA0B4496B204314C3D50426493EE7D4E87C7400628D5A4230EF9AF1C7AEF2BD6EDF0DCD201FD98BA6BC44F93FD46E248AB1C884B1AC28E43BBA2F112125EA2131F84CB932638B5BB442FBCEAF2B47530E0B1B6C13F00956F4B6E7FA63DA1E26AE4E297940EF3F56B9BA6EC55DA6CF9D7A76D03564640FA87250724F9A26E9DD87E524681909AB0DA10C9767A53075D52C5F98F8772998445DE3C3D78DE3B35ACE025421706F7AAE6B99A8A762D89B925997BB0621A9229371EBCF3C7D896A7553C1CFE03477643103C56A4A3A0168A8EBBE5D69E539E4BC7EFA115DEA52DB0B06AD8D8970182172FF0A111D3A99BDEB6BA48DCEEC3B8F1D98A2841C92E6839E7FD71CA60DF13313BF03CAB7D053526F98F8F632DC1C852DE9BBB94B2AE88BDB6FE665114AAB42428A33DED0B5666EDFE1FF88790E1D9AD55CCE0E98DEAC4F14680740860DE1479D48D475F425117CBDB5AB2C6D8AD04534FB2D7415761BC1B24471414D5CB08D79E33AC671E29455E30E12FF2AE378017214ABD2E8784BB759630131994FB547CEC2FD11F676E11C1C1195647270D1015B0701BD2548E2751CBE9947A50E7513A4BF4CD2414BEB75E45E038B4E28333DB58236CB6ADAD7DCD5BE0D169CE4F79F5175436ADF9EF477AC4A58D10D846798C2B528BDC9CACDDC579E630D7D31496BC0BEF028E269B4A25BC7FCA1AB7F36E112C4A8223C016716FA98ADC35AD2AD0232CF7B06D98828DA6F9E2BFA1142B7722924D287C9011914469CA552B8014BDB4A06482AD9A812B9A4F663AB3C46DDEC13BB2735766514436878E9133D27CFB7DBF569DC1021F5E4FF721E7CACA057F40E6C00C9E445D606704A9CF49F37D98BC7955A163196B07A21A568A643B3062B37FA42A2FB20FB9E340E85B97963971F97B34CC9B323E4C4596D6312893C47855DE0232BAD338CC4C0EF59D57DFF1B15B3CA07AB3CB100A2AB9D542C63B0BFAD6D4A5F6FF03760B2B836DDBF955D0CBB810610E200D43D0F3F9A8711ABA08D29D3A772D3E3A7ECE6B669CB2C1A7D0F3B1C273164D00172F7950E4F174D624BAA6F0F938FE3961444B63C2C7E7520F246DE4EFE5E47EC52CFF0417B584E2CA9CBF8058341ECF24BB74C165938FD4AC118384E8356C837592648D50E20E0B5484561DF8637F6B73F79F6A1A2B0E878D7D5F0EE7F7A6D341E9B6BAC6A1D039AF1CE87431A6FD923A9F82703A0C3378368C15658FAD872472DA193D5EBD1F04D6C19AC9C319A66A658A4C574DAC687872F0D8236A71A1CB7AF82CB5F905B2DF6508E02CE2F0CBE76E0CDCCDE4169D05FA137224C398DF307F58E2A38621A17E4E7E07E21C3A4EDACFAC351B3CD3405E1BA9C20D5B9854951EC2A7EE94D87653DA5EDDBD301BE0B8E77D3A27AA879DAA00EACC5EC86C4FEFE49306986EE9D37FF43CA0A7CD1A3B19045BE0C8F23474A32AFA122794B58451E6A403523AA2F014A6D285A0A1F35856E3C218BF6030FE43324394F4AD1CA6BC7C7797C0312FF4B4268B5BE4978EA8C60658F213335A32F89DCF733A90D40F72A5270815013127F196C320469A357302875695A6884C70BCD76D436C148E76C133AE05B52AC4DF1755554C0E10965367752682B7EB25822DBD8DFE365F53C6C0992E8A5D3502C2AB205EE6A97DA24A4E245624BF28919D16205660AC91725F2261E4754FA09F0035BA315FF50946BB8736DE98BEFA544E3C2B412851B24D6269B0084F2CB451B09D77187175ADCD8632B77124845580CE8ADB45AD920B8CE99FF909E8884C8157887D7C54C23BE4C2990DD053CF19C3EE107F1295CF766D7474C4E9162592368742AAA21CCA0E96246E15ACDC282EE646B3C1C8B08266BF13C981F7AA09819BDC57002D773C862875AA516BD93420C3A061DE8C4B1102EAA95921512B8E226511D3DB32606A9D79107F4E3DFB978593D406EB4510CE33EF026B96D12466D155F982ED466F9C68C612664EA0DC65E3762ACBD160992AE9DB6513520A880C6207825EF98FAFAE37BEA4187BD2020EF4FB2A52070B23EA7E252D192F2BFAB5649F1B518E38D8ADC0FA78BAF2ABEB7BBF939B6ED36C666F5C8EE95810B76ACB8DD61D3C38EA3A88C75AA33F8DBB3A49EE813C59205752C8D76910145ED92EE9C2FED1884FCF353187FF0CB92C57D5E4B24DFB3C4F9D0BC5E298063A3E38C818143C3EDB2390AEC7EA8A9C1F7593A47692A4ED28C825AFF73C907044660254E42266B89C6AAEC330476F8E5FF47CC466D91F172C70B05E9142385B64E90B712793568FD607D7045359AF7CE791CC915BF8CD70C620E8BC29E6929F6AC0597A8CFB2D90597A643761C1E9AC1D2474CCF270A373F7B20E9C5ABADFCFCF009DE96DC41173090223C8949120B5E1598CA6AAA0457AFA8B73947E7D23540FE80015CB49B02946CDA39B0F8D686FDF6C6FE65521A300020927D97E8A64B4F7413B6EA67D6EAFDC22C915B28915761FA58E54104A92221648CABCC4DB19935CB3001973BD8852183829267C6ABBDFA2A725BEFDC2226E1A923CF6A0F17C9D73FAD4C1ACE116972411CFD8B8F10E7C29E1F20BE9EF6A78BC5400DCCAA72CAEF22841CFFAD98D91ED33B1FE9BAB0B61E81A38960184FF9AA04C4B96CEDDF84085AAE2953A1652B2ED124D71C54E8FC43834618CFA3D1A7BE6D9C440CF94D8A33210D685BB0BCFF6F4F5FF45FE00515D84331E17FDEE96A3FFB0AA5BFEE4BA012F8449CE8BE46D44876D3FEBB2EA94A7B3DDDB0940B2B42ADFEC0AA7BBD9E273519B899B2E9F4099FF9850D4B2F4F0EB2F37FDD56601480BDAA7B261A26B095AFDEE68E3B0E849F39E1A5E592BD4B949C18F45B6C74E4F7D0CDD2CFFEAA0E2B68CA175443AEC05CBF00346491312EDA4519324CEB0EC589D33AE9BDB35167C3314E5544C5BDDA5635075DF86A16CCF00CF4D808EB6D90FB597250CEDF267DBC71EF69E2F86D23C9C7EF4A6DECA48FFE2A939F108BF04968DEF558921DC24A20EC7C5482C2B2CDF9ED0A99A869CE030356717DC307572CCC956136464EB7543E0FAEC09AA5908554AE7B09BD40A2CB7482F17D497A2FECA7AA57D60A20ED33B30DD84C2C69AE717BC615F4CD7C390D357A6E548673BF3BEB447E76EFBF3A95C67D6DFB1E8018970EF176A7AE638E90E2837259C693B179C9550F38CF686A15A951B1CD52C311A230DA3A70C6659F24BDCF97646F6EDE966EF25C8C90A3293104B66EBADF186BFC762E2D0FFDD3A2FB6C5D6E73D86576B17BD7441F363F8BB4DD0D11C811F892AE3C80F3469130518766D6E8FEE9064D9099AC116B4EF2B0EC4C7B6BAFBB4BF0F862DC789C471B436A9611F490230F292B0D8E996A03C8363A9EB203E6471B09FD273AC878134B4054C3A652C45E9688EB2607B1EFBD1B49F1795353CDC5F05A497A0E86922D5FEE02F0A2943081211733C0C5ED681A1557D8281406FA3908C549175BE4914C9F0A75F8F9EF2E293BB0823DD814059515D69962C0DF1CF1F446E8FD31945F15BD72C19DC77009D1403AAF63A1C651070D55A5EB5E0A98E81C4C2A87531F89EDEF1D78324001AC428CCDC46F6C78DEE65C4630B262A85A0233708A3D1AE16FD5C51912CE521BEA750DAAA1BE19738C397AE03AE7C92B9C5F596ED12071055110AA322A23AA20F841D907367BD377F28AB924973DE45425DDC7657E7F22C43572985788EED02139CA903BF4209F583EA96F1F55A1D70E60F05D591D54B3ECF86C17A65F6A8F3243094E924339FB7BB88750BD1183590773B18F9E437F512E2814DF4ADABDB343754F3162C1514BD92DAEFA69F62860C6E181EDB769D0282DC2F1AF0DC93C62E2DA9ECB2237C7077A1296C5B3ECE592D9A8ADF72898ABFE2FE2D452BBF02690CC01ED8C447C035E61366D4E3A5D33E00E6622B1AAE347D8F84E343A2B532A7FBF49447B9FA6DF35FA0DAD42CA091E736B8AE98AF5171A5B2E36F612A82976CBA37C07A1C843F666881DCA648941A5E5C407CBA33D1C39F19442C80BC94B705999EFBBC579C66C135D0D388381752CB2B3CBBF1C6A4EB731C9C33D7E64B319034765D3CA45C9BC116D10C34C5D4D19F627138A77C60EEC5825337046C20EE6E1CD51E4F6D549F59FDD48C25C8DD1C32414CA7C7A737AC038933E5DAA1D78AE7A59DFB7BAE4EFA9A5A7D7A248781D7439DC4D5A4105A1AEE1AFBB03BAB1E480305354871F78FBA8F7AC10943DADC455380F5ADCF2763BB07931CAFA4B46CD23BB6C65DF5E0E6E40E7AE559307A2973AF04A2B2F4A0361777EC71D4212737916A097CCE070F33792AE73D943D7AEBB55AB0A963C4D11AB678C5F811B924201F0D175F144F04B148EFF1AA2FC9E08712DF48039122C7336AC7EE73C698C3CA8BEDF5205FF70B63901A21818BE59FD88324BD19AD6E662DCB9D3E7B3FAD689DEBCFC4976E76BE92C02BB4FA67AA9E8D22EB5B5B6A8D6CC4E9DB7402C858936C21B2EB68F8A20A6D7F915A0CD8F97AABC677DF86A2FC50E004F660C312E2DF9CF23894484C905ED941D3C6FFD426C9B0ACBBA4E634032AC680F049638C2CCEDA4A2E07BD49C643D2015E656270775C82A3B15DA877F164A6A9D7FD372E7753FF8673322F9C6F337B9B33391C0D1A2E509655C97A25CF0CE6B07334BA684A0ED59843A6534EC31B3C64EED4B4B36D005C9F8C1F0A2D30C52AC272E81C0DCC3FF441F3683294DFD8AA94D53D3BACB1C9627416E41E5246951C6FEFB9F1E5FB8FB38CD1FA7CBEC2ABB01A83F6F20098893F4937B591A5B649027FC698E41FE72DA8AB7C88694E050A2F5AC2BD4B3C54F35D46841B17778EFE8E656BA1698C7AE547928C1CE494A2DDC5B7A110F7ADA124FEF591CB963FE0163022B82A8B1F2EA39D3FCDC1DE1F0069EF47B413EF6DA732FFCD0C1A945EEC14F2CDA4318B5C51202672324FAD91A7F0D2139DFA7FD6813B2CAAE80EA15376622C225189D70599C63D0A6BA56BE56E789D3B69DF51FB38B53497FD25AB1C13C6D82B55D6D4AB87DB7444B20C51124FB1C12AB5C04237F95D13722476999C6E4C30F94892BE8805CDE70C3E11BF9B51E9684AD66FF34DAB72EEE624E3C6137C17D62DD2464AA861C92807F3F8D91D4AB7CF77CD70CB8A64E4BC7CA05BFE2640969604F97176A5DDA043F31AA5AA383FC46EF1138BC1B53F2A31E80DDA1E53B5DB4A03D596E2D377EAA0653FDA62E43008C43A8EAD107BDF3BAFD24E2A57AB5B7D2CCA8610038D7471DCA3572A613EB454124231896D42C74B771C7A60F2CCF93FFFC16E1E66C34CB6D97D275932EF44CD92CC65BC30B1C7B4B62CDE86A6AB342D61EB725DAAA07349CB013084ECE121865ECEF967D982A711ED3CA891E1C8ED61D3AB1A5F4FF76CF3F196CEC304852454AD1A06DE244F214CFBBB413EDDF8EF398E34DEEBD4A58ABC742EAE77708849DA842B4D050E8246929E939A402B9E6486E10F0E53D04A9C4356A08F3D8F52A9B37D743E93DF456DC6DCC87165588317786E10084005FAD84F528328484C11E6F937B9FAE8122C512C526809333C6B129E7E27F4DA66EA1907390465827DD031D061675BF7611BA09FB3A0477C74E2C52C2049B829D5AF689D1946132B78F0841B7585059EBF30CBDE598C98D1C4EB509C6957D68AE34959242497740A31A2E374E03F0620873E85ED7D05F605A0729DA67CB38EB85A6529E95F243BD35D301B7E6E4E3FB930ACBA48CD7AC12B94EFD24F0C2FAE97AD1101852F852F5F65730B350C177EBE1FC2A4D7770A577D867B5A4C5B7040BC6FEC75A5242CD501CCC57B03FD7552D8F0E754F3D8D4FF7414C5126D6C4097FED27DD408D86952DB743AA7461108C1AABE06AFE43ED5293249D86E7E7033D71B1E8A270B205AA84E148B2E22DA9D1D1CC5931C70198FC823FD0BEC5D5C66761B1556D96736BD6AFF1000293DD630C816497C060E34D1539AE990D2E3C84AA60A68DD3609DF51C731CDF9EA3F6BA280A21E3F576B026AABE542D234C81B0C5E8D112F69411FBF6DD7C4DE91F4D11D21AF181F4870430D2E3CA68C0300F7636028BABE21AD19DD51966062433CB79BB9A75EE6EA5A485DC4C60C0A0DBE65E72AAF30033FC76C3EC9DD80A16D3E4D2495B2E6DC618FB7ECC2627BE11755B014018D9D9548FDF17D5F86BE20E8ABF8E8853CC9070E7BF0BDBAF095379BCD37E9D45EE2F7C2E6108C111B61D18D99754DEA8C8CEDF55572D21D8E55979119E20D66EE423EC3F8891088E3B3C9C7F4893B3FFA813C2E30AA446EC01FDA0396A7232DE035DB9A97A9D00A3B506D23FBC02FA83369393A66FF0EBE48EBECB92291205A13549DD06C2DC62AAE7E44CF313EEA7EECD9E52B2F8D493EA47E4D3B0FC991473AB78B385CF83E55497D70602CCECFFFC018F678873F91E8CC93ED7077CBEC66FD546A216EEA1A62C7A23EC58C9F0A835579F014D995BA80D280788C532328CF93B5F7C63B892B64C20CF795868456BF00F7394EDB3304A91DA23504B48BF7910013CA2FFF0CEB4C648FCE3B03C538BDA2C1AE7491B96B2AC8005F9A0E8D65A752166DD22B9DBAA5AE897CBA24CF5BAF64C64269D85718EE4FF5DFE0964A56015B274AEFCD8D962718C30C9DF1E1C5A8A7565257E9ECFA393F45EF92FC6DFCE864F56C54383F409F35FCF481C3FA2AF9DCDF68F874435B3177B1849C7FE22E195DE0BC161701476D06D28B8FC2E25EAF6E77FE4DBAE4DB2C3DD1E05C6AE53B18F2E469E16AE46B5AA5B5EE4BF82FE779B1E2FF2DE500D99BDD6C64842C99874F3DB304BF8807E9E34855E3E7C1B7375AA639C5BB076B579697CB90680EC80D39FDFAD09CB9363251086222E09F41AA07B2A8610E7457257312D4BA7BDF9EFF161E6C308D7C199EAC3292B5D46324CBC8405A97FAF941C9692969CF7A5BD6C448CA671711F1E2F257F35BAC59C0B861ACA52ACB4315E11DD8B98A2E744D54FDD82C0FE78EF498FFD5C25A67D84473613FDC4C687CB38EB437E2A52916CF5E577DEA5886AAF155524F171FBC713308D0EFBBB6D3189403DA234A7CD0C96BC7B373A37A36DF8E205544F7558AE9452959431B57F30537E4EC89C90B958AFE366E3F5A039618881B0A0750E79008AF0441E3FB8BDF0EADF78C5217FC335D4BBC0A1C26EAD379AC3CB5E1994FC724C94B22FBB8CE8F116F9D48D59F21C378AE4579826F6CE9BBC230A7E781FC6E0E01AB42C2418677BEA34CD1628F80939F082C8809BC3F0BF45AD0A19FA1CD32038E01A9EFE73B493911FE09C8D21CE68FE5E9002EB7691D30099A35AF6B8D367FB02A5AF51B74F03FB1AF29D5C66FB72BDA5AD707C1BB35AB6C867B4D423DE1951800BA52F4B855073A8443A25CA227017072DD5F1A428CD2C8326567C933838E8E4C6D31F602A6419DBEA1AB932D91686204B24D3D64BCD'
			},
		]
	},
]
